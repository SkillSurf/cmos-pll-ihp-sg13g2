** T2_VCO_INVERTER flat netlist
*.PININFO VPWR:B VGND:B A:I Y:O VPB:B VNB:B
*--------BEGIN_XM2->SG13_LV_PMOS
XM2 Y A VPWR VPB  SG13_LV_PMOS W=1U L=0.13U NG=1 M=1
*--------END___XM2->SG13_LV_PMOS
*--------BEGIN_XM1->SG13_LV_NMOS
XM1 Y A VGND VNB  SG13_LV_NMOS W=0.5U L=0.13U NG=1 M=1
*--------END___XM1->SG13_LV_NMOS
.end
