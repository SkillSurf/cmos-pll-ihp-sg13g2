** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_and2.sch
.subckt t2_and2 VDD VSS inA out inB
*.PININFO VSS:B inA:I inB:I out:O VDD:B
x1 VDD inA inB net1 VSS t2_nand2
x2 VDD net1 net1 out VSS t2_nand2
.ends

* expanding   symbol:  t2_nand2.sym # of pins=5
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand2.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand2.sch
.subckt t2_nand2 VDD inA inB out VSS
*.PININFO VSS:B inA:I inB:I out:O VDD:B
M1 out inA VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M2 out inB VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M3 out inB net1 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M4 net1 inA VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends

