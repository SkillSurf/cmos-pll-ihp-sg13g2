** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_freq_divider.sch
.subckt t2_freq_divider VDD VSS clk_in en lmt0 lmt1 lmt2 lmt3 clk_out
*.PININFO VSS:B lmt0:I VDD:B clk_out:O lmt1:I lmt2:I lmt3:I clk_in:I en:I
x1 VDD VSS net2 net5 net1 cout0 t2_ha
x2 VDD VSS net1 clk_b div_rst net2 net3 t2_dff_1
x3 VDD VSS net2 lmt0 neq0 t2_xor2
* noconn #net3
x4 VDD VSS net5 net4 t2_tie
* noconn #net4
* noconn clk_out
x5 VDD VSS net6 div_rst net8 clk_out net6 t2_dff_1
x7 VDD VSS net8 net7 t2_tie
* noconn #net7
x8 VDD VSS net10 cout0 net9 cout1 t2_ha
x9 VDD VSS net9 clk_b div_rst net10 net11 t2_dff_1
x10 VDD VSS net10 lmt1 neq1 t2_xor2
* noconn #net11
x11 VDD VSS net13 cout1 net12 cout2 t2_ha
x12 VDD VSS net12 clk_b div_rst net13 net14 t2_dff_1
x13 VDD VSS net13 lmt2 neq2 t2_xor2
* noconn #net14
x14 VDD VSS net16 cout2 net15 net17 t2_ha
x15 VDD VSS net15 clk_b div_rst net16 net18 t2_dff_1
x16 VDD VSS net16 lmt3 neq3 t2_xor2
* noconn #net18
* noconn #net17
x17 VDD VSS neq0 neq1 neq2 neq3 div_rst t2_or4
x6 VDD clk_in en clk_b VSS t2_nand2
.ends

* expanding   symbol:  t2_ha.sym # of pins=6
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_ha.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_ha.sch
.subckt t2_ha VDD VSS inA inB sum cout
*.PININFO VSS:B inA:I inB:I sum:O VDD:B cout:O
x1 VDD VSS inA inB sum t2_xor2
x2 VDD VSS inA cout inB t2_and2
.ends


* expanding   symbol:  t2_dff_1.sym # of pins=7
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_dff_1.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_dff_1.sch
.subckt t2_dff_1 VDD VSS D CLK RST Q QN
*.PININFO VSS:B D:I RST:I Q:O VDD:B QN:O CLK:I
x3 VDD net1 QN Q VSS t2_nand2
x4 VDD VSS Q net2 RST QN t2_nand3
x1 VDD VSS net4 net5 RST net1 t2_nand3
x2 VDD VSS net1 net5 net3 net2 t2_nand3
x6 VDD net3 net1 net4 VSS t2_nand2
x5 VDD VSS net2 D RST net3 t2_nand3
x7 VDD CLK net5 VSS t2_inverter
.ends


* expanding   symbol:  t2_xor2.sym # of pins=5
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_xor2.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_xor2.sch
.subckt t2_xor2 VDD VSS inA inB out
*.PININFO VSS:B inA:I inB:I out:O VDD:B
x1 VDD inA inB net1 VSS t2_nand2
x2 VDD inA net1 net3 VSS t2_nand2
x3 VDD net1 inB net2 VSS t2_nand2
x4 VDD net3 net2 out VSS t2_nand2
.ends


* expanding   symbol:  t2_tie.sym # of pins=4
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_tie.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_tie.sch
.subckt t2_tie VDD VSS outHI outLO
*.PININFO VSS:B outLO:O VDD:B outHI:O
M1 outHI net1 VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M2 net1 net1 VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M3 net2 net2 VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M4 outLO net2 VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  t2_or4.sym # of pins=7
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_or4.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_or4.sch
.subckt t2_or4 VDD VSS inA inB inC inD out
*.PININFO VSS:B inD:I out:O VDD:B inA:I inB:I inC:I
x1 VDD VSS inA inB net2 t2_or2
x2 VDD VSS inC inD net1 t2_or2
x3 VDD VSS net2 net1 out t2_or2
.ends


* expanding   symbol:  t2_nand2.sym # of pins=5
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand2.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand2.sch
.subckt t2_nand2 VDD inA inB out VSS
*.PININFO VSS:B inA:I inB:I out:O VDD:B
M1 out inA VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M2 out inB VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M3 out inB net1 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M4 net1 inA VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  t2_and2.sym # of pins=5
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_and2.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_and2.sch
.subckt t2_and2 VDD VSS inA out inB
*.PININFO VSS:B inA:I inB:I out:O VDD:B
x1 VDD inA inB net1 VSS t2_nand2
x2 VDD net1 net1 out VSS t2_nand2
.ends


* expanding   symbol:  t2_nand3.sym # of pins=6
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand3.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand3.sch
.subckt t2_nand3 VDD VSS inA inB inC out
*.PININFO VSS:B inA:I inC:I out:O VDD:B inB:I
M1 out inB VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M2 out inC VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M3 out inC net1 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M4 net1 inB net2 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M5 net2 inA VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M0 out inA VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  t2_inverter.sym # of pins=4
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_inverter.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_inverter.sch
.subckt t2_inverter VP A Y VN
*.PININFO VP:B VN:B A:I Y:O
M2 Y A VP VP sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M1 Y A VN VN sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  t2_or2.sym # of pins=5
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_or2.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_or2.sch
.subckt t2_or2 VDD VSS inA inB out
*.PININFO VSS:B inA:I inB:I out:O VDD:B
x2 VDD inA inA net2 VSS t2_nand2
x3 VDD inB inB net1 VSS t2_nand2
x4 VDD net2 net1 out VSS t2_nand2
.ends

