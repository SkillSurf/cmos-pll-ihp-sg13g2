* NGSPICE file created from pll_3bitDiv.ext - technology: ihp-sg13g2

.subckt pll_3bitDiv CLK_IN CLK_OUT Y0 Y2 Y1 VDD VSS nEN X1 X2 X0
X0 PFD_0.VDD a_53968_20434# a_53899_20488# PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X1 PFD_0.VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_61488_20220# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X2 a_62119_20605# a_61691_20534# a_61394_20220# PFD_0.VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X3 a_52924_22885# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X4 a_53065_20179# a_53738_20514# a_53702_20612# PFD_0.VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=43.05f ps=0.625u w=0.42u l=0.13u
X5 a_62119_22361# 3bit_freq_divider_1.dff_nclk_0.nCLK PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1533p pd=1.57u as=0.11785p ps=1.025u w=0.42u l=0.13u
X6 PFD_0.VSS a_53152_43159# cap_cmim l=6.99u w=6.99u
X7 PFD_0.VDD a_52950_22157# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q PFD_0.VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X8 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X9 PFD_0.VSS 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_61061_23234# PFD_0.VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.1216p ps=1.02u w=0.64u l=0.13u
X10 a_62879_24125# a_61887_24046# a_62654_23727# PFD_0.VDD sg13_lv_pmos ad=43.05f pd=0.625u as=0.17695p ps=1.56u w=0.42u l=0.13u
X11 a_53022_43738# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X12 PFD_0.VSS a_55345_24897# 3bit_freq_divider_0.freq_div_cell_0.Cin PFD_0.VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X13 a_64383_23434# a_64383_23628# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X14 PFD_0.VDD a_53774_21934# a_53738_22270# PFD_0.VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X15 a_55485_23233# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.1331p ps=1.12u w=0.64u l=0.13u
X16 a_64383_23300# a_64383_23628# a_64424_22200# PFD_0.VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X17 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.53658n ps=1.60669m w=1.5u l=0.65u
X18 PFD_0.VDD a_53022_43738# a_57084_43159# PFD_0.VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X19 PFD_0.VDD a_51648_21103# 3bit_freq_divider_0.dff_nclk_0.nCLK PFD_0.VDD sg13_lv_pmos ad=0.3822p pd=1.84u as=0.3808p ps=2.92u w=1.12u l=0.13u
X20 a_64383_23434# a_64383_23628# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X21 a_54627_42591# 11Stage_vco_new_0.vctl PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X22 a_59799_40285# a_58520_43159# a_58515_40413# PFD_0.VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X23 a_61972_23244# 3bit_freq_divider_1.freq_div_cell_0.Cin PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X24 a_54494_43159# a_53152_43159# a_54627_42591# PFD_0.VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X25 a_54427_40283# a_54489_40413# a_53147_40413# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X26 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D a_54504_23771# PFD_0.VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X27 a_53774_20178# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X28 a_54504_20259# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D a_55086_20219# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X29 charge_pump_0.bias_n charge_pump_0.bias_n PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.34p pd=2.68u as=0.34p ps=2.68u w=1u l=1u
X30 PFD_0.VSS 3bit_freq_divider_0.freq_div_cell_0.Cout a_54434_21392# PFD_0.VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X31 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_63463_23728# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.14505p ps=1.15u w=0.74u l=0.13u
X32 a_47954_28913# PFD_0.VCO_CLK a_48909_28913# PFD_0.VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X33 a_54898_21129# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_54434_21392# PFD_0.VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X34 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X35 a_51693_23426# 3bit_freq_divider_0.dff_nclk_0.nRST PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1533p pd=1.57u as=0.11785p ps=1.025u w=0.42u l=0.13u
X36 PFD_0.VSS a_54489_40413# cap_cmim l=6.99u w=6.99u
X37 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.dff_nclk_0.nCLK PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X38 PFD_0.UP a_47777_29803# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.1632p pd=1.64u as=0.1632p ps=1.64u w=0.48u l=0.15u
X39 PFD_0.VDD a_62654_23727# a_62900_23691# PFD_0.VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=79.8f ps=0.8u w=0.42u l=0.13u
X40 a_54504_23771# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D a_55086_23731# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X41 a_60967_23234# 3bit_freq_divider_1.freq_div_cell_0.Cin PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.2856p ps=2.36u w=0.84u l=0.13u
X42 a_54602_23243# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D PFD_0.VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X43 a_54898_24641# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_54434_24904# PFD_0.VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X44 PFD_0.VDD 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_60967_21478# PFD_0.VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.1596p ps=1.22u w=0.84u l=0.13u
X45 a_62221_24117# a_61691_24046# a_62119_24117# PFD_0.VDD sg13_lv_pmos ad=51.45f pd=0.665u as=79.8f ps=0.8u w=0.42u l=0.13u
X46 a_58426_43159# a_57178_43159# a_58520_43159# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X47 a_62246_20260# a_61887_20534# a_62119_20605# PFD_0.VSS sg13_lv_nmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X48 a_52074_23051# a_51684_22692# a_51693_23426# PFD_0.VSS sg13_lv_nmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X49 a_54504_22015# 3bit_freq_divider_0.dff_nclk_0.nCLK PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X50 PFD_0.VDD a_55345_23141# 3bit_freq_divider_0.freq_div_cell_0.Cout PFD_0.VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X51 a_64464_23130# a_64419_23326# a_64464_23052# PFD_0.VSS sg13_lv_nmos ad=48.3f pd=0.65u as=54.6f ps=0.68u w=0.42u l=0.13u
X52 PFD_0.VSS a_63255_21488# 3bit_freq_divider_1.sg13g2_or3_1_0.A PFD_0.VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X53 a_61675_22886# 3bit_freq_divider_1.freq_div_cell_0.Cin PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X54 PFD_0.VDD a_53022_43738# a_53085_40283# PFD_0.VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X55 a_53968_20434# a_53738_20514# a_54324_20259# PFD_0.VSS sg13_lv_nmos ad=79.8f pd=0.8u as=54.6f ps=0.68u w=0.42u l=0.13u
X56 PFD_0.VSS 3bit_freq_divider_0.sg13g2_or3_1_0.B a_51648_21103# PFD_0.VSS sg13_lv_nmos ad=0.1045p pd=0.93u as=0.198p ps=1.27u w=0.55u l=0.13u
X57 PFD_0.VDD 3bit_freq_divider_0.EN charge_pump_0.bias_p PFD_0.VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X58 a_55345_23141# 3bit_freq_divider_0.freq_div_cell_0.Cin a_55485_23233# PFD_0.VSS sg13_lv_nmos ad=0.2176p pd=1.96u as=0.1216p ps=1.02u w=0.64u l=0.13u
X59 charge_pump_0.bias_n charge_pump_0.bias_p a_55862_56737# PFD_0.VDD sg13_lv_pmos ad=0.68p pd=4.68u as=0.38p ps=2.38u w=2u l=1u
X60 a_53152_43159# a_52944_43077# a_53058_43159# PFD_0.VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X61 PFD_0.VDD a_53022_43738# a_55769_40283# PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X62 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI a_60584_24580# a_60385_24558# PFD_0.VDD sg13_lv_pmos ad=0.3927p pd=2.99u as=0.4657p ps=2.54u w=1.155u l=0.13u
X63 a_54324_20259# a_53899_20488# a_54252_20259# PFD_0.VSS sg13_lv_nmos ad=54.6f pd=0.68u as=48.3f ps=0.65u w=0.42u l=0.13u
X64 a_62270_24055# a_62119_24117# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X65 a_62324_22016# a_62270_22299# a_62246_22016# PFD_0.VSS sg13_lv_nmos ad=48.3f pd=0.65u as=54.6f ps=0.68u w=0.42u l=0.13u
X66 PFD_0.VDD 3bit_freq_divider_0.A2 a_52924_21129# PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X67 3bit_freq_divider_0.CLK_IN a_59614_43129# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X68 a_52944_43077# a_53147_40413# a_53085_40283# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X69 PFD_0.VSS a_53774_21934# a_53738_22270# PFD_0.VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X70 a_46749_30782# PFD_0.Ref_CLK a_45579_29803# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.15u
X71 a_54400_43159# a_53152_43159# a_54494_43159# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X72 3bit_freq_divider_1.freq_div_cell_0.Cin a_60967_24990# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.1918p ps=1.5u w=1.12u l=0.13u
X73 a_55742_43159# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X74 a_53968_23946# a_53738_24026# a_54324_23771# PFD_0.VSS sg13_lv_nmos ad=79.8f pd=0.8u as=54.6f ps=0.68u w=0.42u l=0.13u
X75 a_63038_20215# 3bit_freq_divider_1.dff_nclk_0.nCLK PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=47.25f pd=0.645u as=90.3f ps=0.85u w=0.42u l=0.13u
X76 a_62900_20179# a_62654_20215# a_63038_20215# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=47.25f ps=0.645u w=0.42u l=0.13u
X77 3bit_freq_divider_0.sg13g2_or3_1_0.C a_52886_24904# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X78 PFD_0.VDD a_53022_43738# a_57111_40283# PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X79 a_48909_28913# PFD_0.VCO_CLK a_47954_28913# PFD_0.VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=68.39999f ps=0.74u w=0.36u l=0.15u
X80 a_54324_23771# a_53899_24000# a_54252_23771# PFD_0.VSS sg13_lv_nmos ad=54.6f pd=0.68u as=48.3f ps=0.65u w=0.42u l=0.13u
X81 PFD_0.VSS 11Stage_vco_new_0.vctl a_58454_40850# PFD_0.VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X82 a_58453_40283# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X83 a_53899_22244# a_53774_21934# a_53065_21935# PFD_0.VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.17695p ps=1.56u w=1u l=0.13u
X84 PFD_0.VDD 3bit_freq_divider_0.A0 a_52924_24641# PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X85 PFD_0.VDD a_64384_21091# 3bit_freq_divider_1.dff_nclk_0.nCLK PFD_0.VDD sg13_lv_pmos ad=0.3822p pd=1.84u as=0.3808p ps=2.92u w=1.12u l=0.13u
X86 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_61972_23244# PFD_0.VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X87 PFD_0.VDD 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI a_61878_24642# PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X88 3bit_freq_divider_1.sg13g2_or3_1_0.B a_63255_23244# a_63426_22886# PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X89 PFD_0.VSS 11Stage_vco_new_0.vctl a_53022_43738# PFD_0.VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X90 a_51729_23026# a_51631_22774# a_51693_23426# PFD_0.VDD sg13_lv_pmos ad=51.45f pd=0.665u as=79.8f ps=0.8u w=0.42u l=0.13u
X91 a_57084_43159# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X92 a_61887_20534# a_61691_20534# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X93 a_54400_43159# a_53152_43159# a_54494_43159# PFD_0.VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X94 a_62119_22361# a_61691_22290# a_61394_21976# PFD_0.VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X95 a_52950_23913# a_53065_23691# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.2016p ps=1.5u w=0.84u l=0.13u
X96 a_54504_20259# a_53738_20514# a_53968_20434# PFD_0.VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X97 a_62119_24117# 3bit_freq_divider_1.dff_nclk_0.nCLK PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1533p pd=1.57u as=0.11785p ps=1.025u w=0.42u l=0.13u
X98 PFD_0.VCO_CLK PFD_0.VCO_CLK a_46817_27899# PFD_0.VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X99 PFD_0.VDD 3bit_freq_divider_0.CLK_IN 3bit_freq_divider_1.sg13g2_nand2_1_0.Y PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X100 PFD_0.VSS 3bit_freq_divider_0.CLK_IN cap_cmim l=6.99u w=6.99u
X101 PFD_0.VDD a_62900_21935# a_62879_22369# PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=43.05f ps=0.625u w=0.42u l=0.13u
X102 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X103 a_53350_21129# 3bit_freq_divider_0.A2 a_52886_21392# PFD_0.VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X104 a_58454_40850# a_58515_40413# a_57173_40413# PFD_0.VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X105 PFD_0.VSS 3bit_freq_divider_0.EN a_56055_21027# PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=66.6f ps=0.92u w=0.74u l=0.13u
X106 PFD_0.VDD a_62654_23727# a_63463_23728# PFD_0.VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.2856p ps=2.36u w=0.84u l=0.13u
X107 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X108 a_55742_43159# a_54494_43159# a_55836_43159# PFD_0.VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X109 a_62654_21971# a_61887_22290# a_62270_22299# PFD_0.VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=0.19397p ps=1.29u w=0.64u l=0.13u
X110 PFD_0.VSS a_62900_20179# a_62848_20215# PFD_0.VSS sg13_lv_nmos ad=90.3f pd=0.85u as=54.6f ps=0.68u w=0.42u l=0.13u
X111 PFD_0.VSS 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X112 a_61394_23732# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X113 a_62848_20215# a_61691_20534# a_62654_20215# PFD_0.VSS sg13_lv_nmos ad=54.6f pd=0.68u as=0.2017p ps=1.48u w=0.42u l=0.13u
X114 PFD_0.VSS a_58515_40413# cap_cmim l=6.99u w=6.99u
X115 a_53774_21934# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X116 a_53054_23243# 3bit_freq_divider_0.A1 3bit_freq_divider_0.sg13g2_or3_1_0.B PFD_0.VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X117 a_53350_24641# 3bit_freq_divider_0.A0 a_52886_24904# PFD_0.VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X118 PFD_0.VDD a_53022_43738# a_58426_43159# PFD_0.VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X119 a_56038_24617# a_55941_24882# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI PFD_0.VDD sg13_lv_pmos ad=0.4657p pd=2.54u as=0.3927p ps=2.99u w=1.155u l=0.13u
X120 PFD_0.VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53445_20214# PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X121 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X122 a_57112_40850# 11Stage_vco_new_0.vctl PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X123 a_60584_24580# a_60385_24717# a_60479_25023# PFD_0.VSS sg13_lv_nmos ad=0.27427p pd=2.28u as=0.2307p ps=1.615u w=0.795u l=0.13u
X124 PFD_0.VSS a_61707_21488# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D PFD_0.VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X125 a_63255_25000# 3bit_freq_divider_1.A0 a_63223_24642# PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X126 PFD_0.VDD a_51648_24041# a_51685_23725# PFD_0.VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=79.8f ps=0.8u w=0.42u l=0.13u
X127 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_63463_20216# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2016p ps=1.5u w=1.12u l=0.13u
X128 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D a_54434_21392# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X129 PFD_0.VSS 3bit_freq_divider_1.A0 a_63255_25000# PFD_0.VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X130 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X131 a_48909_28913# PFD_0.VCO_CLK a_47954_28913# PFD_0.VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=0.1224p ps=1.4u w=0.36u l=0.15u
X132 PFD_0.VDD a_62270_20543# a_62221_20605# PFD_0.VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=51.45f ps=0.665u w=0.42u l=0.13u
X133 a_62246_22016# a_61887_22290# a_62119_22361# PFD_0.VSS sg13_lv_nmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X134 PFD_0.VDD 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_63426_21130# PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X135 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_0.Cout a_54898_21129# PFD_0.VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X136 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X137 a_64362_24865# a_64459_24995# a_64731_24890# PFD_0.VDD sg13_lv_pmos ad=0.2442p pd=2.06u as=0.4657p ps=2.54u w=0.66u l=0.13u
X138 a_55831_40413# a_57173_40413# a_57112_40850# PFD_0.VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X139 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X140 a_47777_29803# a_46749_30782# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=0.1224p ps=1.4u w=0.36u l=0.15u
X141 a_55086_21975# 3bit_freq_divider_0.dff_nclk_0.nCLK PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X142 PFD_0.VDD 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_54898_24641# PFD_0.VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X143 a_53445_21970# a_53065_21935# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.2163p ps=1.55u w=0.42u l=0.13u
X144 PFD_0.VSS 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_52886_23148# PFD_0.VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X145 a_64384_21091# 3bit_freq_divider_1.sg13g2_or3_1_0.A PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.198p pd=1.27u as=0.13395p ps=1.12u w=0.55u l=0.13u
X146 a_63255_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X147 a_54494_43159# a_53152_43159# a_54400_43159# PFD_0.VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X148 a_63426_24642# 3bit_freq_divider_1.A0 PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X149 a_62270_20543# a_62119_20605# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.1825p ps=1.325u w=0.64u l=0.13u
X150 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X151 PFD_0.VSS 11Stage_vco_new_0.vctl a_58653_42591# PFD_0.VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X152 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ a_62654_21971# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2775p pd=2.23u as=0.2516p ps=2.16u w=0.74u l=0.13u
X153 a_58653_42591# a_57178_43159# a_58520_43159# PFD_0.VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X154 PFD_0.VDD a_64383_23889# a_64384_24445# PFD_0.VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.2856p ps=2.36u w=0.84u l=0.13u
X155 a_51708_21299# 3bit_freq_divider_0.sg13g2_or3_1_0.A PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.22p pd=1.44u as=0.3822p ps=1.84u w=1u l=0.13u
X156 PFD_0.VSS 3bit_freq_divider_0.dff_nclk_0.nRST a_52074_23129# PFD_0.VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=48.3f ps=0.65u w=0.42u l=0.13u
X157 a_53147_40413# a_54489_40413# a_54427_40283# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X158 PFD_0.VDD 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X159 PFD_0.VSS a_57178_43159# cap_cmim l=6.99u w=6.99u
X160 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.51p pd=3.68u as=0 ps=0 w=1.5u l=0.65u
X161 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X162 PFD_0.VSS a_53147_40413# cap_cmim l=6.99u w=6.99u
X163 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X164 a_62879_20613# a_61887_20534# a_62654_20215# PFD_0.VDD sg13_lv_pmos ad=43.05f pd=0.625u as=0.17695p ps=1.56u w=0.42u l=0.13u
X165 a_61887_22290# a_61691_22290# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X166 PFD_0.VSS a_52950_22157# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q PFD_0.VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.2516p ps=2.16u w=0.74u l=0.13u
X167 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X168 a_63520_25000# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X169 a_53702_24124# a_53445_23726# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=43.05f pd=0.625u as=79.8f ps=0.8u w=0.42u l=0.13u
X170 a_61707_25000# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X171 PFD_0.VDD 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_22290# PFD_0.VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X172 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_54472_21129# PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X173 PFD_0.VSS 3bit_freq_divider_0.freq_div_cell_0.Cin a_54602_23243# PFD_0.VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X174 PFD_0.VSS a_51648_24041# a_51648_24438# PFD_0.VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.187p ps=1.78u w=0.55u l=0.13u
X175 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X176 a_53147_40413# a_54489_40413# a_54427_40283# PFD_0.VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X177 a_62270_20543# a_62119_20605# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X178 a_51648_21103# 3bit_freq_divider_0.sg13g2_or3_1_0.C a_51708_21413# PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1275p ps=1.255u w=1u l=0.13u
X179 PFD_0.VDD 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_51631_22774# PFD_0.VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X180 PFD_0.VSS 11Stage_vco_new_0.vctl a_53086_40850# PFD_0.VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X181 a_59800_40852# 11Stage_vco_new_0.vctl PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X182 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X183 a_53085_40283# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X184 a_62654_23727# a_61887_24046# a_62270_24055# PFD_0.VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=0.19397p ps=1.29u w=0.64u l=0.13u
X185 3bit_freq_divider_0.EN sg13g2_inv_1_0.A PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X186 PFD_0.VDD a_58734_56203# a_58734_56203# PFD_0.VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X187 PFD_0.VDD a_64383_23706# a_64817_23685# PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=43.05f ps=0.625u w=0.42u l=0.13u
X188 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_54472_24641# PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X189 PFD_0.VSS 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X190 a_55862_56737# PFD_0.VDD rhigh l=12u w=1u
X191 PFD_0.VDD a_46817_27899# a_45658_27900# PFD_0.VDD sg13_lv_pmos ad=0.1224p pd=1.4u as=68.39999f ps=0.74u w=0.36u l=0.15u
X192 3bit_freq_divider_1.sg13g2_or3_1_0.B 3bit_freq_divider_1.A1 a_63520_23244# PFD_0.VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X193 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X194 a_54489_40413# a_55831_40413# a_55769_40283# PFD_0.VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X195 a_57084_43159# a_55836_43159# a_57178_43159# PFD_0.VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X196 a_63223_24642# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X197 a_58520_43159# a_57178_43159# a_58426_43159# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X198 a_58515_40413# a_58520_43159# a_59800_40852# PFD_0.VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X199 PFD_0.VDD a_62654_20215# a_62900_20179# PFD_0.VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=79.8f ps=0.8u w=0.42u l=0.13u
X200 a_53086_40850# a_53147_40413# a_52944_43077# PFD_0.VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X201 a_64424_22294# 3bit_freq_divider_1.dff_nclk_0.D a_64424_22200# PFD_0.VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X202 a_61488_23732# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D a_61394_23732# PFD_0.VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X203 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X204 a_61061_21478# 3bit_freq_divider_1.freq_div_cell_0.Cout a_60967_21478# PFD_0.VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.2176p ps=1.96u w=0.64u l=0.13u
X205 PFD_0.VSS 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_51631_22774# PFD_0.VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X206 a_62221_20605# a_61691_20534# a_62119_20605# PFD_0.VDD sg13_lv_pmos ad=51.45f pd=0.665u as=79.8f ps=0.8u w=0.42u l=0.13u
X207 PFD_0.VSS a_53968_22190# a_53899_22244# PFD_0.VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=0.19397p ps=1.29u w=0.64u l=0.13u
X208 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X209 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.CLK_IN a_60531_21028# PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=66.6f ps=0.92u w=0.74u l=0.13u
X210 PFD_0.VDD a_53022_43738# a_54427_40283# PFD_0.VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X211 PFD_0.VSS a_55345_21385# 3bit_freq_divider_0.freq_div_cell_1.Cout PFD_0.VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X212 a_59097_54704# 3bit_freq_divider_0.EN PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X213 PFD_0.VSS a_55831_40413# cap_cmim l=6.99u w=6.99u
X214 a_52114_22293# 3bit_freq_divider_0.dff_nclk_0.D a_51684_22284# PFD_0.VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X215 a_51693_23075# a_51693_23426# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X216 PFD_0.VDD a_64383_23889# a_64383_23706# PFD_0.VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=79.8f ps=0.8u w=0.42u l=0.13u
X217 a_61061_24990# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI a_60967_24990# PFD_0.VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.2176p ps=1.96u w=0.64u l=0.13u
X218 a_54472_21129# 3bit_freq_divider_0.freq_div_cell_0.Cout PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X219 a_61887_22290# a_61691_22290# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X220 PFD_0.VDD a_53022_43738# a_53058_43159# PFD_0.VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X221 3bit_freq_divider_0.CLK_IN a_59614_43129# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X222 a_61878_24642# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X223 PFD_0.VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_61488_21976# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X224 a_54400_43159# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X225 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_63463_20216# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.14505p ps=1.15u w=0.74u l=0.13u
X226 a_54434_23148# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X227 PFD_0.VDD a_53022_43738# a_55769_40283# PFD_0.VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X228 3bit_freq_divider_0.dff_nclk_0.D a_51648_24041# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.7616p pd=3.6u as=0.2163p ps=1.55u w=1.12u l=0.13u
X229 3bit_freq_divider_1.freq_div_cell_0.Cout a_60967_23234# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1331p ps=1.12u w=0.74u l=0.13u
X230 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X231 a_54472_24641# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X232 a_55485_24989# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.1331p ps=1.12u w=0.64u l=0.13u
X233 PFD_0.VCO_CLK a_51648_24438# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.14505p ps=1.15u w=0.74u l=0.13u
X234 a_62900_21935# 3bit_freq_divider_1.dff_nclk_0.nCLK PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X235 a_53774_21934# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X236 a_55742_43159# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X237 a_53899_22244# a_53738_22270# a_53065_21935# PFD_0.VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.2017p ps=1.48u w=0.64u l=0.13u
X238 a_64383_23889# a_64383_23628# a_64419_23326# PFD_0.VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=0.19p ps=1.38u w=1u l=0.13u
X239 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ a_62654_23727# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2775p pd=2.23u as=0.2516p ps=2.16u w=0.74u l=0.13u
X240 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.dff_nclk_0.nCLK PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X241 a_58426_43159# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X242 PFD_0.VSS 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_53054_23243# PFD_0.VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X243 PFD_0.VSS 3bit_freq_divider_1.A2 a_63255_21488# PFD_0.VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X244 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X245 PFD_0.VDD a_59614_43129# 3bit_freq_divider_0.CLK_IN PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X246 a_52950_20401# a_53065_20179# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.2016p ps=1.5u w=0.84u l=0.13u
X247 a_62119_20605# 3bit_freq_divider_1.dff_nclk_0.nCLK PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1533p pd=1.57u as=0.11785p ps=1.025u w=0.42u l=0.13u
X248 a_60531_21028# 3bit_freq_divider_0.EN PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=66.6f pd=0.92u as=0.2516p ps=2.16u w=0.74u l=0.13u
X249 PFD_0.VDD a_52950_20401# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q PFD_0.VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X250 a_47777_29803# a_46749_30782# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1224p pd=1.4u as=68.39999f ps=0.74u w=0.36u l=0.15u
X251 PFD_0.VSS a_52950_23913# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q PFD_0.VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.2516p ps=2.16u w=0.74u l=0.13u
X252 a_51693_23075# a_51693_23426# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.1825p ps=1.325u w=0.64u l=0.13u
X253 PFD_0.VDD 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_24046# PFD_0.VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X254 a_54602_24999# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D PFD_0.VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X255 a_53065_21935# a_53738_22270# a_53702_22368# PFD_0.VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=43.05f ps=0.625u w=0.42u l=0.13u
X256 PFD_0.VSS 11Stage_vco_new_0.vctl a_53285_42591# PFD_0.VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X257 PFD_0.VDD a_62654_20215# a_63463_20216# PFD_0.VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.2856p ps=2.36u w=0.84u l=0.13u
X258 a_53285_42591# a_52944_43077# a_53152_43159# PFD_0.VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X259 PFD_0.VDD 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_60967_23234# PFD_0.VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.1596p ps=1.22u w=0.84u l=0.13u
X260 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D a_61707_25000# a_61878_24642# PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X261 3bit_freq_divider_1.freq_div_cell_1.Cout a_60967_21478# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.1918p ps=1.5u w=1.12u l=0.13u
X262 a_54842_49733# a_54357_49278# charge_pump_0.vout PFD_0.VDD sg13_lv_pmos ad=55.5f pd=0.74u as=0.1005p ps=1.34u w=0.15u l=0.13u
X263 PFD_0.VSS a_54494_43159# cap_cmim l=6.99u w=6.99u
X264 a_61707_25000# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_61675_24642# PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X265 a_61394_20220# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X266 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D a_54504_22015# PFD_0.VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X267 a_55345_23141# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.1918p ps=1.5u w=0.84u l=0.13u
X268 charge_pump_0.bias_n sg13g2_inv_1_0.A PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X269 a_53022_43738# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X270 PFD_0.VSS 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_61707_25000# PFD_0.VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X271 3bit_freq_divider_0.sg13g2_or3_1_0.A a_52886_21392# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X272 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X273 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X274 a_54427_40283# a_54489_40413# a_53147_40413# PFD_0.VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X275 a_54252_20259# 3bit_freq_divider_0.dff_nclk_0.nCLK PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=48.3f pd=0.65u as=0.1825p ps=1.325u w=0.42u l=0.13u
X276 a_55345_24897# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_55485_24989# PFD_0.VSS sg13_lv_nmos ad=0.2176p pd=1.96u as=0.1216p ps=1.02u w=0.64u l=0.13u
X277 3bit_freq_divider_1.CLK_OUT a_64384_24445# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.14505p ps=1.15u w=0.74u l=0.13u
X278 a_54504_20259# a_53774_20178# a_53968_20434# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X279 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X280 PFD_0.VSS a_51685_23725# a_52119_23653# PFD_0.VSS sg13_lv_nmos ad=90.3f pd=0.85u as=54.6f ps=0.68u w=0.42u l=0.13u
X281 PFD_0.VDD 3bit_freq_divider_1.freq_div_cell_0.Cout a_61878_21130# PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X282 a_52950_22157# a_53065_21935# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.187p pd=1.78u as=0.14505p ps=1.15u w=0.55u l=0.13u
X283 a_55969_42591# 11Stage_vco_new_0.vctl PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X284 a_54427_40283# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X285 a_55836_43159# a_54494_43159# a_55969_42591# PFD_0.VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X286 a_55770_40850# 11Stage_vco_new_0.vctl PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X287 a_62654_23727# a_61691_24046# a_62270_24055# PFD_0.VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=0.19p ps=1.38u w=1u l=0.13u
X288 a_64714_21414# 3bit_freq_divider_1.sg13g2_or3_1_0.B a_64714_21300# PFD_0.VDD sg13_lv_pmos ad=0.1275p pd=1.255u as=0.22p ps=1.44u w=1u l=0.13u
X289 PFD_0.VDD a_51648_24041# a_51648_24438# PFD_0.VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.2856p ps=2.36u w=0.84u l=0.13u
X290 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X291 a_52924_21129# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X292 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X293 a_55769_40283# a_55831_40413# a_54489_40413# PFD_0.VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X294 a_54252_23771# 3bit_freq_divider_0.dff_nclk_0.nCLK PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=48.3f pd=0.65u as=0.1825p ps=1.325u w=0.42u l=0.13u
X295 PFD_0.VSS a_62654_21971# a_63463_21972# PFD_0.VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.187p ps=1.78u w=0.55u l=0.13u
X296 PFD_0.VDD a_45658_27900# PFD_0.DOWN PFD_0.VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X297 3bit_freq_divider_1.dff_nclk_0.D a_64383_23889# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.7616p pd=3.6u as=0.2163p ps=1.55u w=1.12u l=0.13u
X298 a_45658_27900# a_46817_27899# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=68.39999f pd=0.74u as=0.1224p ps=1.4u w=0.36u l=0.15u
X299 PFD_0.VSS 3bit_freq_divider_0.dff_nclk_0.nCLK a_53539_21970# PFD_0.VSS sg13_lv_nmos ad=90.3f pd=0.85u as=47.25f ps=0.645u w=0.42u l=0.13u
X300 a_53539_21970# a_53065_21935# a_53445_21970# PFD_0.VSS sg13_lv_nmos ad=47.25f pd=0.645u as=0.1428p ps=1.52u w=0.42u l=0.13u
X301 PFD_0.VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53968_22190# PFD_0.VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=0.1533p ps=1.57u w=0.42u l=0.13u
X302 a_54504_23771# a_53774_23690# a_53968_23946# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X303 PFD_0.VSS a_53968_23946# a_53899_24000# PFD_0.VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=0.19397p ps=1.29u w=0.64u l=0.13u
X304 a_52924_22885# a_52886_23148# 3bit_freq_divider_0.sg13g2_or3_1_0.B PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X305 a_52886_23148# 3bit_freq_divider_0.A1 PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X306 a_58453_40283# a_58515_40413# a_57173_40413# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X307 a_63520_21488# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X308 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ a_62654_23727# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.7616p pd=3.6u as=0.2163p ps=1.55u w=1.12u l=0.13u
X309 a_64731_24890# a_64398_24796# 3bit_freq_divider_1.dff_nclk_0.nRST PFD_0.VDD sg13_lv_pmos ad=0.4657p pd=2.54u as=0.3927p ps=2.99u w=1.155u l=0.13u
X310 a_61707_21488# 3bit_freq_divider_1.freq_div_cell_0.Cout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X311 a_54427_40283# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X312 PFD_0.VDD a_53968_22190# a_53899_22244# PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X313 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X314 a_52924_24641# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X315 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X316 a_54489_40413# a_55831_40413# a_55770_40850# PFD_0.VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X317 PFD_0.VDD a_52950_23913# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q PFD_0.VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X318 a_61887_24046# a_61691_24046# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X319 charge_pump_0.vout 11Stage_vco_new_0.vctl rhigh l=0.96u w=0.6u
X320 PFD_0.VDD a_53065_21935# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ PFD_0.VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=0.7616p ps=3.6u w=1.12u l=0.13u
X321 a_53152_43159# a_52944_43077# a_53058_43159# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X322 PFD_0.VDD a_51685_23725# a_51721_23684# PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=43.05f ps=0.625u w=0.42u l=0.13u
X323 PFD_0.VDD a_53774_23690# a_53738_24026# PFD_0.VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X324 a_55836_43159# a_54494_43159# a_55742_43159# PFD_0.VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X325 a_55769_40283# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X326 a_56013_24979# a_56137_24678# a_56038_24617# PFD_0.VDD sg13_lv_pmos ad=0.2442p pd=2.06u as=0.4657p ps=2.54u w=0.66u l=0.13u
X327 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_0.Cin a_55345_23141# PFD_0.VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.1596p ps=1.22u w=0.84u l=0.13u
X328 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X329 a_48909_28913# PFD_0.Ref_CLK PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=0.1224p ps=1.4u w=0.36u l=0.15u
X330 a_64464_23052# a_64383_23434# a_64383_23300# PFD_0.VSS sg13_lv_nmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X331 a_56055_21027# 3bit_freq_divider_0.CLK_IN 3bit_freq_divider_0.sg13g2_nand2_1_0.Y PFD_0.VSS sg13_lv_nmos ad=66.6f pd=0.92u as=0.2516p ps=2.16u w=0.74u l=0.13u
X332 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X333 a_61972_25000# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X334 a_63255_21488# 3bit_freq_divider_1.A2 a_63223_21130# PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X335 a_51648_21103# 3bit_freq_divider_0.sg13g2_or3_1_0.C PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.187p pd=1.78u as=0.1045p ps=0.93u w=0.55u l=0.13u
X336 a_53899_24000# a_53738_24026# a_53065_23691# PFD_0.VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.2017p ps=1.48u w=0.64u l=0.13u
X337 PFD_0.VSS 3bit_freq_divider_0.freq_div_cell_0.Cin a_54434_23148# PFD_0.VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X338 charge_pump_0.vout PFD_0.DOWN a_54747_49259# PFD_0.VSS sg13_lv_nmos ad=0.408p pd=3.08u as=0.207p ps=1.545u w=1.2u l=0.13u
X339 a_52119_23843# 3bit_freq_divider_0.dff_nclk_0.nRST PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=47.25f pd=0.645u as=90.3f ps=0.85u w=0.42u l=0.13u
X340 PFD_0.UP a_47777_29803# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X341 a_53054_24999# 3bit_freq_divider_0.A0 3bit_freq_divider_0.sg13g2_or3_1_0.C PFD_0.VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X342 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X343 a_57178_43159# a_55836_43159# a_57084_43159# PFD_0.VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X344 PFD_0.VDD a_55345_21385# 3bit_freq_divider_0.freq_div_cell_1.Cout PFD_0.VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X345 PFD_0.VDD 3bit_freq_divider_1.dff_nclk_0.nCLK a_61394_23732# PFD_0.VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X346 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X347 a_57084_43159# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X348 a_53065_21935# a_53774_21934# a_53722_21970# PFD_0.VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=54.6f ps=0.68u w=0.42u l=0.13u
X349 a_53968_22190# a_53774_21934# a_54352_22360# PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=51.45f ps=0.665u w=0.42u l=0.13u
X350 a_53702_20612# a_53445_20214# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=43.05f pd=0.625u as=79.8f ps=0.8u w=0.42u l=0.13u
X351 PFD_0.VDD a_53022_43738# a_58426_43159# PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X352 PFD_0.VSS 11Stage_vco_new_0.vctl a_59800_40852# PFD_0.VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X353 a_59799_40285# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X354 a_60967_24990# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.2856p ps=2.36u w=0.84u l=0.13u
X355 PFD_0.VDD a_53022_43738# a_53085_40283# PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X356 a_53722_21970# a_53445_21970# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=54.6f pd=0.68u as=90.3f ps=0.85u w=0.42u l=0.13u
X357 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X358 PFD_0.VSS 11Stage_vco_new_0.vctl a_54428_40850# PFD_0.VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X359 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X360 PFD_0.VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_62324_23772# PFD_0.VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=48.3f ps=0.65u w=0.42u l=0.13u
X361 PFD_0.VDD a_55345_24897# 3bit_freq_divider_0.freq_div_cell_0.Cin PFD_0.VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X362 PFD_0.VSS a_63255_23244# 3bit_freq_divider_1.sg13g2_or3_1_0.B PFD_0.VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X363 a_61675_24642# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X364 a_53058_43159# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X365 PFD_0.VDD 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_63426_22886# PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X366 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.CLK_IN PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X367 a_53968_22190# a_53738_22270# a_54324_22015# PFD_0.VSS sg13_lv_nmos ad=79.8f pd=0.8u as=54.6f ps=0.68u w=0.42u l=0.13u
X368 a_63426_21130# 3bit_freq_divider_1.A2 PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X369 a_61394_21976# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X370 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X371 PFD_0.VSS a_59600_42432# 3bit_freq_divider_0.CLK_IN PFD_0.VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X372 a_54324_22015# a_53899_22244# a_54252_22015# PFD_0.VSS sg13_lv_nmos ad=54.6f pd=0.68u as=48.3f ps=0.65u w=0.42u l=0.13u
X373 a_59800_40852# a_58520_43159# a_58515_40413# PFD_0.VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X374 a_58734_56203# a_58536_54976# a_58536_54976# PFD_0.VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X375 a_54428_40850# a_54489_40413# a_53147_40413# PFD_0.VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X376 a_52950_23913# a_53065_23691# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.187p pd=1.78u as=0.14505p ps=1.15u w=0.55u l=0.13u
X377 a_64383_23300# a_64383_23434# a_64424_22200# PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X378 PFD_0.VSS 3bit_freq_divider_1.sg13g2_or3_1_0.B a_64384_21091# PFD_0.VSS sg13_lv_nmos ad=0.1045p pd=0.93u as=0.198p ps=1.27u w=0.55u l=0.13u
X379 PFD_0.VSS 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_52886_24904# PFD_0.VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X380 PFD_0.VDD 3bit_freq_divider_0.dff_nclk_0.nRST a_51684_22284# PFD_0.VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X381 PFD_0.VDD charge_pump_0.bias_p charge_pump_0.bias_p PFD_0.VDD sg13_lv_pmos ad=0.68p pd=4.68u as=0.68p ps=4.68u w=2u l=1u
X382 a_64459_24995# a_64459_24995# a_64338_24910# PFD_0.VSS sg13_lv_nmos ad=0.102p pd=1.28u as=0.2307p ps=1.615u w=0.3u l=0.13u
X383 PFD_0.VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53445_21970# PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X384 PFD_0.VDD PFD_0.UP a_54357_49278# PFD_0.VDD sg13_lv_pmos ad=0.102p pd=1.28u as=0.102p ps=1.28u w=0.3u l=0.13u
X385 PFD_0.VSS a_62654_23727# a_63463_23728# PFD_0.VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.187p ps=1.78u w=0.55u l=0.13u
X386 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X387 a_53899_24000# a_53774_23690# a_53065_23691# PFD_0.VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.17695p ps=1.56u w=1u l=0.13u
X388 PFD_0.VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53968_23946# PFD_0.VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=0.1533p ps=1.57u w=0.42u l=0.13u
X389 a_53539_23726# a_53065_23691# a_53445_23726# PFD_0.VSS sg13_lv_nmos ad=47.25f pd=0.645u as=0.1428p ps=1.52u w=0.42u l=0.13u
X390 PFD_0.VSS 3bit_freq_divider_0.dff_nclk_0.nCLK a_53539_23726# PFD_0.VSS sg13_lv_nmos ad=90.3f pd=0.85u as=47.25f ps=0.645u w=0.42u l=0.13u
X391 a_57311_42591# 11Stage_vco_new_0.vctl PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X392 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_61972_25000# PFD_0.VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X393 3bit_freq_divider_1.sg13g2_or3_1_0.C a_63255_25000# a_63426_24642# PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X394 a_57178_43159# a_55836_43159# a_57311_42591# PFD_0.VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X395 a_45579_29803# PFD_0.Ref_CLK a_45451_28860# PFD_0.VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=68.39999f ps=0.74u w=0.36u l=0.15u
X396 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_63463_21972# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2016p ps=1.5u w=1.12u l=0.13u
X397 PFD_0.VSS 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_24046# PFD_0.VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X398 PFD_0.VSS 3bit_freq_divider_0.CLK_IN cap_cmim l=6.99u w=6.99u
X399 PFD_0.VDD 3bit_freq_divider_1.dff_nclk_0.nRST a_64424_22200# PFD_0.VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X400 PFD_0.VDD a_64419_23326# a_64809_23027# PFD_0.VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=51.45f ps=0.665u w=0.42u l=0.13u
X401 a_64338_24910# a_64362_24865# a_64398_24796# PFD_0.VSS sg13_lv_nmos ad=0.2307p pd=1.615u as=0.27427p ps=2.28u w=0.795u l=0.13u
X402 a_62654_20215# a_61887_20534# a_62270_20543# PFD_0.VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=0.19397p ps=1.29u w=0.64u l=0.13u
X403 PFD_0.DOWN a_45658_27900# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=60.8f pd=0.7u as=60.8f ps=0.7u w=0.32u l=0.15u
X404 a_54472_22885# a_54434_23148# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X405 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_53350_22885# PFD_0.VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X406 PFD_0.VSS 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X407 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X408 a_51648_24041# a_51684_22692# a_51693_23075# PFD_0.VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=0.19397p ps=1.29u w=0.64u l=0.13u
X409 PFD_0.VDD a_62900_23691# a_62879_24125# PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=43.05f ps=0.625u w=0.42u l=0.13u
X410 PFD_0.VSS 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_61707_21488# PFD_0.VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X411 a_45579_29803# PFD_0.Ref_CLK a_45451_28860# PFD_0.VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X412 PFD_0.VSS 3bit_freq_divider_1.dff_nclk_0.nRST a_64424_22294# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X413 a_45579_29803# PFD_0.Ref_CLK PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X414 PFD_0.VSS 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_54602_24999# PFD_0.VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X415 a_63223_21130# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X416 a_58515_40413# a_58520_43159# a_59799_40285# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X417 a_53085_40283# a_53147_40413# a_52944_43077# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X418 a_58515_40413# a_58520_43159# a_59799_40285# PFD_0.VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X419 a_61488_20220# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D a_61394_20220# PFD_0.VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X420 a_62654_20215# a_61691_20534# a_62270_20543# PFD_0.VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=0.19p ps=1.38u w=1u l=0.13u
X421 a_54494_43159# a_53152_43159# a_54400_43159# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X422 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X423 a_55742_43159# a_54494_43159# a_55836_43159# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X424 a_46817_27899# PFD_0.VCO_CLK a_47954_28913# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.15u
X425 PFD_0.VSS 3bit_freq_divider_0.dff_nclk_0.nRST a_52114_22293# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X426 PFD_0.VSS a_53065_21935# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.2775p ps=2.23u w=0.74u l=0.13u
X427 PFD_0.VDD a_53022_43738# a_58453_40283# PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X428 a_54352_22360# a_53899_22244# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=51.45f pd=0.665u as=0.11785p ps=1.025u w=0.42u l=0.13u
X429 PFD_0.VSS a_61707_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D PFD_0.VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X430 PFD_0.VSS a_58520_43159# cap_cmim l=6.99u w=6.99u
X431 a_54357_49278# PFD_0.UP PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.1005p pd=1.34u as=0.1005p ps=1.34u w=0.15u l=0.13u
X432 a_53968_23946# a_53774_23690# a_54352_24116# PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=51.45f ps=0.665u w=0.42u l=0.13u
X433 PFD_0.VDD 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X434 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0 ps=0 w=0.5u l=0.65u
X435 a_53065_23691# a_53774_23690# a_53722_23726# PFD_0.VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=54.6f ps=0.68u w=0.42u l=0.13u
X436 a_61878_21130# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X437 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D a_54434_23148# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X438 PFD_0.VDD 3bit_freq_divider_0.EN a_58536_54976# PFD_0.VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X439 a_57084_43159# a_55836_43159# a_57178_43159# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X440 PFD_0.VDD 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_20534# PFD_0.VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X441 a_53722_23726# a_53445_23726# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=54.6f pd=0.68u as=90.3f ps=0.85u w=0.42u l=0.13u
X442 a_55086_20219# 3bit_freq_divider_0.dff_nclk_0.nCLK PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X443 a_58520_43159# a_57178_43159# a_58426_43159# PFD_0.VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X444 PFD_0.UP a_47777_29803# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X445 a_62879_22369# a_61887_22290# a_62654_21971# PFD_0.VDD sg13_lv_pmos ad=43.05f pd=0.625u as=0.17695p ps=1.56u w=0.42u l=0.13u
X446 PFD_0.VDD a_47777_29803# PFD_0.UP PFD_0.VDD sg13_lv_pmos ad=60.8f pd=0.7u as=60.8f ps=0.7u w=0.32u l=0.15u
X447 PFD_0.VSS 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_61061_21478# PFD_0.VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.1216p ps=1.02u w=0.64u l=0.13u
X448 a_51600_24907# a_51622_24863# 3bit_freq_divider_0.dff_nclk_0.nRST PFD_0.VDD sg13_lv_pmos ad=0.4657p pd=2.54u as=0.3927p ps=2.99u w=1.155u l=0.13u
X449 PFD_0.VSS 3bit_freq_divider_1.dff_nclk_0.nRST a_64464_23130# PFD_0.VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=48.3f ps=0.65u w=0.42u l=0.13u
X450 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0 ps=0 w=0.5u l=0.65u
X451 PFD_0.VDD a_46749_30782# a_47777_29803# PFD_0.VDD sg13_lv_pmos ad=68.39999f pd=0.74u as=0.1224p ps=1.4u w=0.36u l=0.15u
X452 a_55485_21477# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.1331p ps=1.12u w=0.64u l=0.13u
X453 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X454 PFD_0.VSS 11Stage_vco_new_0.vctl a_55969_42591# PFD_0.VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X455 a_55969_42591# a_54494_43159# a_55836_43159# PFD_0.VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X456 PFD_0.VSS 11Stage_vco_new_0.vctl a_55770_40850# PFD_0.VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X457 a_53022_43738# 11Stage_vco_new_0.vctl PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X458 a_55769_40283# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X459 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ a_62654_20215# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2775p pd=2.23u as=0.2516p ps=2.16u w=0.74u l=0.13u
X460 a_55086_23731# 3bit_freq_divider_0.dff_nclk_0.nCLK PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X461 PFD_0.VSS 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_61061_24990# PFD_0.VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.1216p ps=1.02u w=0.64u l=0.13u
X462 PFD_0.VSS a_64383_23706# a_64419_23654# PFD_0.VSS sg13_lv_nmos ad=90.3f pd=0.85u as=54.6f ps=0.68u w=0.42u l=0.13u
X463 a_61972_21488# 3bit_freq_divider_1.freq_div_cell_0.Cout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X464 PFD_0.VDD a_53022_43738# a_53058_43159# PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X465 PFD_0.VSS 11Stage_vco_new_0.vctl PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.1005p pd=1.34u as=0 ps=0 w=0.15u l=0.13u
X466 a_54434_24904# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X467 a_53445_23726# a_53065_23691# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.2163p ps=1.55u w=0.42u l=0.13u
X468 a_54400_43159# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X469 a_51684_22692# a_51631_22774# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X470 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X471 a_57111_40283# a_57173_40413# a_55831_40413# PFD_0.VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X472 a_63255_25000# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X473 charge_pump_0.bias_p a_58536_54976# a_59097_54704# PFD_0.VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X474 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X475 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.dff_nclk_0.nCLK PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X476 PFD_0.VSS a_52950_20401# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q PFD_0.VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.2516p ps=2.16u w=0.74u l=0.13u
X477 PFD_0.VSS 11Stage_vco_new_0.vctl a_57112_40850# PFD_0.VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X478 a_62119_22361# a_61887_22290# a_61394_21976# PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X479 a_64383_23706# 3bit_freq_divider_1.dff_nclk_0.nRST PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X480 a_57111_40283# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X481 a_51693_23426# a_51684_22692# a_51684_22284# PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X482 a_58454_40850# 11Stage_vco_new_0.vctl PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X483 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ a_62654_20215# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.7616p pd=3.6u as=0.2163p ps=1.55u w=1.12u l=0.13u
X484 PFD_0.VDD a_62654_21971# a_62900_21935# PFD_0.VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=79.8f ps=0.8u w=0.42u l=0.13u
X485 a_54504_22015# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D a_55086_21975# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X486 a_55770_40850# a_55831_40413# a_54489_40413# PFD_0.VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X487 a_54602_21487# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D PFD_0.VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X488 a_56039_25022# a_56013_24979# a_55941_24882# PFD_0.VSS sg13_lv_nmos ad=0.2307p pd=1.615u as=0.27427p ps=2.28u w=0.795u l=0.13u
X489 a_51685_23725# a_51648_24041# a_52119_23843# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=47.25f ps=0.645u w=0.42u l=0.13u
X490 a_54898_22885# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_54434_23148# PFD_0.VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X491 a_51693_23426# a_51631_22774# a_51684_22284# PFD_0.VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X492 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X493 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D a_61707_21488# a_61878_21130# PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X494 PFD_0.VSS 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_64383_23628# PFD_0.VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X495 PFD_0.VSS 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_53054_24999# PFD_0.VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X496 a_61887_20534# a_61691_20534# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X497 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X498 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X499 a_64714_21300# 3bit_freq_divider_1.sg13g2_or3_1_0.A PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.22p pd=1.44u as=0.3822p ps=1.84u w=1u l=0.13u
X500 a_54504_20259# 3bit_freq_divider_0.dff_nclk_0.nCLK PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X501 a_61707_21488# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_61675_21130# PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X502 PFD_0.VDD 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_64383_23628# PFD_0.VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X503 a_51684_22692# a_51631_22774# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X504 a_57111_40283# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X505 a_57112_40850# a_57173_40413# a_55831_40413# PFD_0.VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X506 PFD_0.VDD a_53774_20178# a_53738_20514# PFD_0.VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X507 PFD_0.VDD a_51693_23075# a_51729_23026# PFD_0.VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=51.45f ps=0.665u w=0.42u l=0.13u
X508 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X509 a_45451_28860# PFD_0.Ref_CLK a_45579_29803# PFD_0.VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X510 a_55345_21385# 3bit_freq_divider_0.freq_div_cell_0.Cout a_55485_21477# PFD_0.VSS sg13_lv_nmos ad=0.2176p pd=1.96u as=0.1216p ps=1.02u w=0.64u l=0.13u
X511 a_57173_40413# a_58515_40413# a_58454_40850# PFD_0.VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X512 charge_pump_0.bias_p charge_pump_0.bias_n a_56742_53480# PFD_0.VSS sg13_lv_nmos ad=0.34p pd=2.68u as=0.34p ps=2.68u w=1u l=1u
X513 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X514 a_62270_22299# a_62119_22361# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X515 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X516 a_64817_23685# a_64383_23434# a_64383_23889# PFD_0.VDD sg13_lv_pmos ad=43.05f pd=0.625u as=0.17695p ps=1.56u w=0.42u l=0.13u
X517 a_51648_24041# a_51631_22774# a_51693_23075# PFD_0.VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=0.19p ps=1.38u w=1u l=0.13u
X518 PFD_0.VDD a_45658_27900# PFD_0.DOWN PFD_0.VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X519 3bit_freq_divider_1.freq_div_cell_0.Cout a_60967_23234# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.1918p ps=1.5u w=1.12u l=0.13u
X520 a_64419_23844# 3bit_freq_divider_1.dff_nclk_0.nRST PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=47.25f pd=0.645u as=90.3f ps=0.85u w=0.42u l=0.13u
X521 3bit_freq_divider_1.sg13g2_or3_1_0.C 3bit_freq_divider_1.A0 a_63520_25000# PFD_0.VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X522 PFD_0.VSS a_64383_23889# a_64384_24445# PFD_0.VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.187p ps=1.78u w=0.55u l=0.13u
X523 a_64384_21091# 3bit_freq_divider_1.sg13g2_or3_1_0.C a_64714_21414# PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1275p ps=1.255u w=1u l=0.13u
X524 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X525 PFD_0.VSS a_53968_20434# a_53899_20488# PFD_0.VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=0.19397p ps=1.29u w=0.64u l=0.13u
X526 a_45451_28860# PFD_0.Ref_CLK a_45579_29803# PFD_0.VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X527 PFD_0.VDD 3bit_freq_divider_1.dff_nclk_0.nCLK a_61394_20220# PFD_0.VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X528 PFD_0.VSS a_53065_23691# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.2775p ps=2.23u w=0.74u l=0.13u
X529 a_53899_20488# a_53774_20178# a_53065_20179# PFD_0.VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.17695p ps=1.56u w=1u l=0.13u
X530 a_52074_23129# a_51693_23075# a_52074_23051# PFD_0.VSS sg13_lv_nmos ad=48.3f pd=0.65u as=54.6f ps=0.68u w=0.42u l=0.13u
X531 a_62324_23772# a_62270_24055# a_62246_23772# PFD_0.VSS sg13_lv_nmos ad=48.3f pd=0.65u as=54.6f ps=0.68u w=0.42u l=0.13u
X532 PFD_0.VDD PFD_0.Ref_CLK a_45579_29803# PFD_0.VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X533 a_54352_24116# a_53899_24000# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=51.45f pd=0.665u as=0.11785p ps=1.025u w=0.42u l=0.13u
X534 PFD_0.VDD 3bit_freq_divider_0.A1 a_52924_22885# PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X535 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_61972_21488# PFD_0.VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X536 PFD_0.VDD 3bit_freq_divider_1.freq_div_cell_0.Cin a_61878_22886# PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X537 PFD_0.VSS a_53774_23690# a_53738_24026# PFD_0.VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X538 a_54489_40413# a_55831_40413# a_55769_40283# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X539 a_61061_23234# 3bit_freq_divider_1.freq_div_cell_0.Cin a_60967_23234# PFD_0.VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.2176p ps=1.96u w=0.64u l=0.13u
X540 a_55862_56737# charge_pump_0.bias_p charge_pump_0.bias_n PFD_0.VDD sg13_lv_pmos ad=0.38p pd=2.38u as=0.68p ps=4.68u w=2u l=1u
X541 a_62900_21935# a_62654_21971# a_63038_21971# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=47.25f ps=0.645u w=0.42u l=0.13u
X542 a_63038_21971# 3bit_freq_divider_1.dff_nclk_0.nCLK PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=47.25f pd=0.645u as=90.3f ps=0.85u w=0.42u l=0.13u
X543 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X544 3bit_freq_divider_0.dff_nclk_0.D a_51648_24041# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2775p pd=2.23u as=0.2516p ps=2.16u w=0.74u l=0.13u
X545 a_51721_24988# a_51721_24988# a_52065_24890# PFD_0.VSS sg13_lv_nmos ad=0.102p pd=1.28u as=0.2307p ps=1.615u w=0.3u l=0.13u
X546 PFD_0.VSS a_55345_23141# 3bit_freq_divider_0.freq_div_cell_0.Cout PFD_0.VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X547 a_52886_24904# 3bit_freq_divider_0.A0 PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X548 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X549 a_55831_40413# a_57173_40413# a_57111_40283# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X550 a_54504_23771# 3bit_freq_divider_0.dff_nclk_0.nCLK PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X551 a_62119_24117# a_61691_24046# a_61394_23732# PFD_0.VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X552 PFD_0.VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_61488_23732# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X553 3bit_freq_divider_0.EN sg13g2_inv_1_0.A PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X554 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X555 a_59799_40285# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X556 a_53899_20488# a_53738_20514# a_53065_20179# PFD_0.VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.2017p ps=1.48u w=0.64u l=0.13u
X557 PFD_0.VSS PFD_0.VCO_CLK a_45451_28860# PFD_0.VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=0.1224p ps=1.4u w=0.36u l=0.15u
X558 PFD_0.VSS a_46817_27899# a_45658_27900# PFD_0.VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=0.1224p ps=1.4u w=0.36u l=0.15u
X559 a_53054_21487# 3bit_freq_divider_0.A2 3bit_freq_divider_0.sg13g2_or3_1_0.A PFD_0.VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X560 a_53350_22885# 3bit_freq_divider_0.A1 a_52886_23148# PFD_0.VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X561 PFD_0.VSS 11Stage_vco_new_0.vctl a_57311_42591# PFD_0.VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X562 a_62900_23691# 3bit_freq_divider_1.dff_nclk_0.nCLK PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X563 a_53774_23690# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X564 a_57311_42591# a_55836_43159# a_57178_43159# PFD_0.VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X565 a_58653_42591# 11Stage_vco_new_0.vctl PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X566 a_55831_40413# a_57173_40413# a_57111_40283# PFD_0.VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X567 a_60967_21478# 3bit_freq_divider_1.freq_div_cell_0.Cout PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.2856p ps=2.36u w=0.84u l=0.13u
X568 PFD_0.VSS a_62900_21935# a_62848_21971# PFD_0.VSS sg13_lv_nmos ad=90.3f pd=0.85u as=54.6f ps=0.68u w=0.42u l=0.13u
X569 a_58426_43159# a_57178_43159# a_58520_43159# PFD_0.VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X570 a_58520_43159# a_57178_43159# a_58653_42591# PFD_0.VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X571 PFD_0.VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53968_20434# PFD_0.VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=0.1533p ps=1.57u w=0.42u l=0.13u
X572 a_62119_24117# a_61887_24046# a_61394_23732# PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X573 a_54747_49259# charge_pump_0.bias_n PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.207p pd=1.545u as=0.408p ps=3.08u w=1.2u l=0.13u
X574 PFD_0.VDD a_53022_43738# a_54400_43159# PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X575 3bit_freq_divider_0.CLK_IN a_59600_42432# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X576 PFD_0.VDD a_53022_43738# a_53022_43738# PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X577 PFD_0.VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_62324_20260# PFD_0.VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=48.3f ps=0.65u w=0.42u l=0.13u
X578 a_62848_21971# a_61691_22290# a_62654_21971# PFD_0.VSS sg13_lv_nmos ad=54.6f pd=0.68u as=0.2017p ps=1.48u w=0.42u l=0.13u
X579 a_63255_23244# 3bit_freq_divider_1.A1 a_63223_22886# PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X580 a_53774_23690# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X581 PFD_0.VSS 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_54434_24904# PFD_0.VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X582 a_60385_24558# a_60385_24947# a_60385_24717# PFD_0.VDD sg13_lv_pmos ad=0.4657p pd=2.54u as=0.2442p ps=2.06u w=0.66u l=0.13u
X583 PFD_0.VSS 3bit_freq_divider_1.A1 a_63255_23244# PFD_0.VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X584 a_58453_40283# a_58515_40413# a_57173_40413# PFD_0.VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X585 a_46749_30782# PFD_0.Ref_CLK PFD_0.Ref_CLK PFD_0.VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X586 a_61675_21130# 3bit_freq_divider_1.freq_div_cell_0.Cout PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X587 a_52119_23653# a_51631_22774# a_51648_24041# PFD_0.VSS sg13_lv_nmos ad=54.6f pd=0.68u as=0.2017p ps=1.48u w=0.42u l=0.13u
X588 a_52950_22157# a_53065_21935# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.2016p ps=1.5u w=0.84u l=0.13u
X589 PFD_0.VCO_CLK a_51648_24438# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2016p ps=1.5u w=1.12u l=0.13u
X590 3bit_freq_divider_1.dff_nclk_0.D a_64383_23889# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2775p pd=2.23u as=0.2516p ps=2.16u w=0.74u l=0.13u
X591 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X592 PFD_0.VDD a_62900_20179# a_62879_20613# PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=43.05f ps=0.625u w=0.42u l=0.13u
X593 a_55345_21385# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.1918p ps=1.5u w=0.84u l=0.13u
X594 PFD_0.VDD a_53065_20179# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ PFD_0.VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=0.7616p ps=3.6u w=1.12u l=0.13u
X595 a_51648_21103# 3bit_freq_divider_0.sg13g2_or3_1_0.A PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.198p pd=1.27u as=0.13395p ps=1.12u w=0.55u l=0.13u
X596 PFD_0.VSS a_51648_21103# 3bit_freq_divider_0.dff_nclk_0.nCLK PFD_0.VSS sg13_lv_nmos ad=0.13395p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X597 a_52944_43077# a_53147_40413# a_53085_40283# PFD_0.VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X598 a_59799_40285# a_58520_43159# a_58515_40413# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X599 a_53065_23691# a_53738_24026# a_53702_24124# PFD_0.VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=43.05f ps=0.625u w=0.42u l=0.13u
X600 a_54504_22015# a_53738_22270# a_53968_22190# PFD_0.VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X601 PFD_0.VDD a_53022_43738# a_54400_43159# PFD_0.VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X602 PFD_0.VDD a_62654_21971# a_63463_21972# PFD_0.VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.2856p ps=2.36u w=0.84u l=0.13u
X603 a_47954_28913# PFD_0.VCO_CLK PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X604 PFD_0.VDD 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_60967_24990# PFD_0.VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.1596p ps=1.22u w=0.84u l=0.13u
X605 a_52950_20401# a_53065_20179# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.187p pd=1.78u as=0.14505p ps=1.15u w=0.55u l=0.13u
X606 a_53086_40850# 11Stage_vco_new_0.vctl PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X607 a_62246_23772# a_61887_24046# a_62119_24117# PFD_0.VSS sg13_lv_nmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X608 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_0.Cin a_54898_22885# PFD_0.VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X609 PFD_0.VDD a_53022_43738# a_57111_40283# PFD_0.VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X610 a_48909_28913# PFD_0.VCO_CLK a_47954_28913# PFD_0.VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X611 PFD_0.VSS 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_52886_21392# PFD_0.VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X612 a_55345_24897# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.1918p ps=1.5u w=0.84u l=0.13u
X613 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X614 a_58453_40283# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X615 3bit_freq_divider_0.sg13g2_or3_1_0.B a_52886_23148# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X616 PFD_0.VSS a_62654_20215# a_63463_20216# PFD_0.VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.187p ps=1.78u w=0.55u l=0.13u
X617 a_63255_21488# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X618 a_54252_22015# 3bit_freq_divider_0.dff_nclk_0.nCLK PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=48.3f pd=0.65u as=0.1825p ps=1.325u w=0.42u l=0.13u
X619 a_63426_22886# 3bit_freq_divider_1.A1 PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X620 PFD_0.VDD a_53022_43738# a_55742_43159# PFD_0.VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X621 a_51685_23725# 3bit_freq_divider_0.dff_nclk_0.nRST PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X622 a_53539_20214# a_53065_20179# a_53445_20214# PFD_0.VSS sg13_lv_nmos ad=47.25f pd=0.645u as=0.1428p ps=1.52u w=0.42u l=0.13u
X623 PFD_0.VSS 3bit_freq_divider_0.dff_nclk_0.nCLK a_53539_20214# PFD_0.VSS sg13_lv_nmos ad=90.3f pd=0.85u as=47.25f ps=0.645u w=0.42u l=0.13u
X624 PFD_0.VDD 3bit_freq_divider_0.EN 3bit_freq_divider_0.sg13g2_nand2_1_0.Y PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X625 a_54504_22015# a_53774_21934# a_53968_22190# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X626 3bit_freq_divider_1.sg13g2_or3_1_0.A a_63255_21488# a_63426_21130# PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X627 a_52924_21129# a_52886_21392# 3bit_freq_divider_0.sg13g2_or3_1_0.A PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X628 PFD_0.VDD 3bit_freq_divider_1.dff_nclk_0.nCLK a_61394_21976# PFD_0.VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X629 a_57178_43159# a_55836_43159# a_57084_43159# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X630 PFD_0.VSS 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_20534# PFD_0.VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X631 a_53968_20434# a_53774_20178# a_54352_20604# PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=51.45f ps=0.665u w=0.42u l=0.13u
X632 a_64419_23326# a_64383_23300# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.1825p ps=1.325u w=0.64u l=0.13u
X633 a_52944_43077# a_53147_40413# a_53086_40850# PFD_0.VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X634 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.EN PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X635 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X636 a_47954_28913# PFD_0.VCO_CLK a_46817_27899# PFD_0.VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.15u
X637 a_62270_22299# a_62119_22361# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.1825p ps=1.325u w=0.64u l=0.13u
X638 a_62900_23691# a_62654_23727# a_63038_23727# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=47.25f ps=0.645u w=0.42u l=0.13u
X639 a_63038_23727# 3bit_freq_divider_1.dff_nclk_0.nCLK PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=47.25f pd=0.645u as=90.3f ps=0.85u w=0.42u l=0.13u
X640 PFD_0.VDD a_53022_43738# a_53022_43738# PFD_0.VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X641 a_52924_24641# a_52886_24904# 3bit_freq_divider_0.sg13g2_or3_1_0.C PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X642 a_56137_24678# a_56137_24678# a_56039_25022# PFD_0.VSS sg13_lv_nmos ad=0.102p pd=1.28u as=0.2307p ps=1.615u w=0.3u l=0.13u
X643 PFD_0.VSS a_52944_43077# cap_cmim l=6.99u w=6.99u
X644 a_45579_29803# PFD_0.Ref_CLK a_45451_28860# PFD_0.VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=0.1224p ps=1.4u w=0.36u l=0.15u
X645 PFD_0.VSS a_45658_27900# PFD_0.DOWN PFD_0.VSS sg13_lv_nmos ad=0.1632p pd=1.64u as=0.1632p ps=1.64u w=0.48u l=0.15u
X646 a_53702_22368# a_53445_21970# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=43.05f pd=0.625u as=79.8f ps=0.8u w=0.42u l=0.13u
X647 a_63520_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X648 a_61707_23244# 3bit_freq_divider_1.freq_div_cell_0.Cin PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X649 PFD_0.VDD a_59614_43129# 3bit_freq_divider_0.CLK_IN PFD_0.VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X650 a_51759_25014# a_51721_24988# a_51600_24907# PFD_0.VDD sg13_lv_pmos ad=0.2442p pd=2.06u as=0.4657p ps=2.54u w=0.66u l=0.13u
X651 PFD_0.VDD a_53968_23946# a_53899_24000# PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X652 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_0.Cout a_55345_21385# PFD_0.VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.1596p ps=1.22u w=0.84u l=0.13u
X653 PFD_0.VSS 3bit_freq_divider_0.freq_div_cell_0.Cout a_54602_21487# PFD_0.VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X654 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X655 a_53058_43159# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X656 PFD_0.VSS a_64384_21091# 3bit_freq_divider_1.dff_nclk_0.nCLK PFD_0.VSS sg13_lv_nmos ad=0.13395p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X657 PFD_0.VDD a_62270_22299# a_62221_22361# PFD_0.VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=51.45f ps=0.665u w=0.42u l=0.13u
X658 PFD_0.VSS 11Stage_vco_new_0.vctl a_54627_42591# PFD_0.VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X659 a_51721_23684# a_51684_22692# a_51648_24041# PFD_0.VDD sg13_lv_pmos ad=43.05f pd=0.625u as=0.17695p ps=1.56u w=0.42u l=0.13u
X660 a_54627_42591# a_53152_43159# a_54494_43159# PFD_0.VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X661 a_51684_22284# 3bit_freq_divider_0.dff_nclk_0.D PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X662 a_61887_24046# a_61691_24046# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X663 PFD_0.VDD a_53065_23691# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ PFD_0.VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=0.7616p ps=3.6u w=1.12u l=0.13u
X664 a_53445_20214# a_53065_20179# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.2163p ps=1.55u w=0.42u l=0.13u
X665 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X666 PFD_0.VDD 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_55345_24897# PFD_0.VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.1596p ps=1.22u w=0.84u l=0.13u
X667 3bit_freq_divider_1.sg13g2_or3_1_0.A 3bit_freq_divider_1.A2 a_63520_21488# PFD_0.VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X668 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_54472_22885# PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X669 3bit_freq_divider_1.CLK_OUT a_64384_24445# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2016p ps=1.5u w=1.12u l=0.13u
X670 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X671 a_53065_20179# a_53774_20178# a_53722_20214# PFD_0.VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=54.6f ps=0.68u w=0.42u l=0.13u
X672 a_64424_22200# 3bit_freq_divider_1.dff_nclk_0.D PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X673 a_63223_22886# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X674 a_61488_21976# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D a_61394_21976# PFD_0.VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X675 PFD_0.VSS a_62900_23691# a_62848_23727# PFD_0.VSS sg13_lv_nmos ad=90.3f pd=0.85u as=54.6f ps=0.68u w=0.42u l=0.13u
X676 a_53722_20214# a_53445_20214# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=54.6f pd=0.68u as=90.3f ps=0.85u w=0.42u l=0.13u
X677 a_64383_23706# a_64383_23889# a_64419_23844# PFD_0.VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=47.25f ps=0.645u w=0.42u l=0.13u
X678 PFD_0.VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_62324_22016# PFD_0.VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=48.3f ps=0.65u w=0.42u l=0.13u
X679 a_62848_23727# a_61691_24046# a_62654_23727# PFD_0.VSS sg13_lv_nmos ad=54.6f pd=0.68u as=0.2017p ps=1.48u w=0.42u l=0.13u
X680 PFD_0.VDD charge_pump_0.bias_p a_54842_49733# PFD_0.VDD sg13_lv_pmos ad=0.1005p pd=1.34u as=55.5f ps=0.74u w=0.15u l=0.13u
X681 PFD_0.VSS a_56887_49467# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X682 a_46817_27899# PFD_0.VCO_CLK PFD_0.VCO_CLK PFD_0.VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X683 a_57173_40413# a_58515_40413# a_58453_40283# PFD_0.VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X684 a_64384_21091# 3bit_freq_divider_1.sg13g2_or3_1_0.C PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.187p pd=1.78u as=0.1045p ps=0.93u w=0.55u l=0.13u
X685 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X686 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.51p pd=3.68u as=0 ps=0 w=1.5u l=0.65u
X687 a_53285_42591# 11Stage_vco_new_0.vctl PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X688 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D a_54434_24904# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X689 a_54504_23771# a_53738_24026# a_53968_23946# PFD_0.VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X690 PFD_0.VSS a_57173_40413# cap_cmim l=6.99u w=6.99u
X691 a_61878_22886# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X692 PFD_0.Ref_CLK PFD_0.Ref_CLK a_46749_30782# PFD_0.VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X693 a_53058_43159# a_52944_43077# a_53152_43159# PFD_0.VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X694 a_53152_43159# a_52944_43077# a_53285_42591# PFD_0.VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X695 a_54434_21392# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X696 PFD_0.VSS a_63255_25000# 3bit_freq_divider_1.sg13g2_or3_1_0.C PFD_0.VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X697 a_47954_28913# PFD_0.VCO_CLK a_48909_28913# PFD_0.VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X698 PFD_0.VDD 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_63426_24642# PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X699 3bit_freq_divider_1.freq_div_cell_1.Cout a_60967_21478# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1331p ps=1.12u w=0.74u l=0.13u
X700 a_53085_40283# a_53147_40413# a_52944_43077# PFD_0.VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X701 a_54472_22885# 3bit_freq_divider_0.freq_div_cell_0.Cin PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X702 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X703 a_64383_23300# 3bit_freq_divider_1.dff_nclk_0.nRST PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.1533p pd=1.57u as=0.11785p ps=1.025u w=0.42u l=0.13u
X704 a_55769_40283# a_55831_40413# a_54489_40413# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X705 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_63463_21972# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.14505p ps=1.15u w=0.74u l=0.13u
X706 a_54428_40850# 11Stage_vco_new_0.vctl PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X707 PFD_0.VDD PFD_0.VCO_CLK a_47954_28913# PFD_0.VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X708 a_54352_20604# a_53899_20488# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=51.45f pd=0.665u as=0.11785p ps=1.025u w=0.42u l=0.13u
X709 charge_pump_0.vout a_56887_49467# rhigh l=0.96u w=0.5u
X710 a_55836_43159# a_54494_43159# a_55742_43159# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X711 PFD_0.VDD a_53022_43738# a_58453_40283# PFD_0.VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X712 3bit_freq_divider_1.freq_div_cell_0.Cin a_60967_24990# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1331p ps=1.12u w=0.74u l=0.13u
X713 PFD_0.VSS 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_53054_21487# PFD_0.VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X714 PFD_0.VSS 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_22290# PFD_0.VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X715 PFD_0.VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53445_23726# PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X716 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X717 a_54472_21129# a_54434_21392# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X718 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_53350_21129# PFD_0.VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X719 a_57111_40283# a_57173_40413# a_55831_40413# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X720 a_52065_24890# a_51759_25014# a_51622_24863# PFD_0.VSS sg13_lv_nmos ad=0.2307p pd=1.615u as=0.27427p ps=2.28u w=0.795u l=0.13u
X721 a_62270_24055# a_62119_24117# PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.1825p ps=1.325u w=0.64u l=0.13u
X722 a_58426_43159# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X723 a_57173_40413# a_58515_40413# a_58453_40283# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X724 PFD_0.VDD a_53022_43738# a_59799_40285# PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X725 a_64383_23889# a_64383_23434# a_64419_23326# PFD_0.VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=0.19397p ps=1.29u w=0.64u l=0.13u
X726 a_53085_40283# a_53022_43738# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X727 PFD_0.VDD a_53022_43738# a_59799_40285# PFD_0.VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X728 a_62221_22361# a_61691_22290# a_62119_22361# PFD_0.VDD sg13_lv_pmos ad=51.45f pd=0.665u as=79.8f ps=0.8u w=0.42u l=0.13u
X729 a_56742_53480# PFD_0.VSS rhigh l=12u w=1u
X730 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_63463_23728# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2016p ps=1.5u w=1.12u l=0.13u
X731 PFD_0.VDD a_53022_43738# a_54427_40283# PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X732 a_53147_40413# a_54489_40413# a_54428_40850# PFD_0.VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X733 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D a_61707_23244# a_61878_22886# PFD_0.VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X734 PFD_0.VDD a_62270_24055# a_62221_24117# PFD_0.VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=51.45f ps=0.665u w=0.42u l=0.13u
X735 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X736 a_54472_24641# a_54434_24904# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D PFD_0.VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X737 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_53350_24641# PFD_0.VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X738 a_53058_43159# a_52944_43077# a_53152_43159# PFD_0.VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X739 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D a_54504_20259# PFD_0.VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X740 a_61707_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_61675_22886# PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X741 a_64419_23326# a_64383_23300# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X742 a_51708_21413# 3bit_freq_divider_0.sg13g2_or3_1_0.B a_51708_21299# PFD_0.VDD sg13_lv_pmos ad=0.1275p pd=1.255u as=0.22p ps=1.44u w=1u l=0.13u
X743 PFD_0.VSS 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_61707_23244# PFD_0.VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X744 PFD_0.VSS a_53065_20179# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ PFD_0.VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.2775p ps=2.23u w=0.74u l=0.13u
X745 a_62324_20260# a_62270_20543# a_62246_20260# PFD_0.VSS sg13_lv_nmos ad=48.3f pd=0.65u as=54.6f ps=0.68u w=0.42u l=0.13u
X746 a_62900_20179# 3bit_freq_divider_1.dff_nclk_0.nCLK PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X747 PFD_0.VSS a_55836_43159# cap_cmim l=6.99u w=6.99u
X748 a_53774_20178# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X749 PFD_0.VSS a_53774_20178# a_53738_20514# PFD_0.VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X750 PFD_0.VDD a_53022_43738# a_55742_43159# PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X751 a_45579_29803# PFD_0.Ref_CLK a_46749_30782# PFD_0.VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.15u
X752 a_62119_20605# a_61887_20534# a_61394_20220# PFD_0.VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X753 a_62654_21971# a_61691_22290# a_62270_22299# PFD_0.VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=0.19p ps=1.38u w=1u l=0.13u
X754 a_60479_25023# a_60385_24947# a_60385_24947# PFD_0.VSS sg13_lv_nmos ad=0.2307p pd=1.615u as=0.102p ps=1.28u w=0.3u l=0.13u
X755 a_64809_23027# a_64383_23628# a_64383_23300# PFD_0.VDD sg13_lv_pmos ad=51.45f pd=0.665u as=79.8f ps=0.8u w=0.42u l=0.13u
X756 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.dff_nclk_0.nCLK PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X757 a_64419_23654# a_64383_23628# a_64383_23889# PFD_0.VSS sg13_lv_nmos ad=54.6f pd=0.68u as=0.2017p ps=1.48u w=0.42u l=0.13u
X758 PFD_0.VSS 11Stage_vco_new_0.vctl PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.1005p pd=1.34u as=0 ps=0 w=0.15u l=0.13u
X759 a_52886_21392# 3bit_freq_divider_0.A2 PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X760 a_58536_54976# charge_pump_0.bias_n PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.34p pd=2.68u as=0.34p ps=2.68u w=1u l=1u
X761 PFD_0.VSS a_61707_25000# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D PFD_0.VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X762 PFD_0.VDD a_53022_43738# a_57084_43159# PFD_0.VDD sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X763 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ a_62654_21971# PFD_0.VDD PFD_0.VDD sg13_lv_pmos ad=0.7616p pd=3.6u as=0.2163p ps=1.55u w=1.12u l=0.13u
X764 PFD_0.VDD 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X765 PFD_0.VSS charge_pump_0.vout PFD_0.VSS PFD_0.VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
C0 a_56828_53480# a_56742_53480# 0.09853f
C1 a_51759_25014# 3bit_freq_divider_0.dff_nclk_0.nRST 0.03098f
C2 a_47777_29803# PFD_0.UP 0.62819f
C3 PFD_0.VDD a_52950_22157# 0.2364f
C4 a_64384_24445# 3bit_freq_divider_1.dff_nclk_0.nRST 0.04054f
C5 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.11142f
C6 3bit_freq_divider_1.A1 m6_17427_2840# 1.19758f
C7 a_53774_21934# a_53738_22270# 0.44698f
C8 a_64383_23434# PFD_0.VDD 0.19308f
C9 3bit_freq_divider_0.dff_nclk_0.nCLK a_53738_24026# 0.18638f
C10 a_63426_24642# 3bit_freq_divider_1.A0 0.01851f
C11 a_63255_23244# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.10223f
C12 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 0.21745f
C13 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_0.Cout 0.42266f
C14 3bit_freq_divider_0.dff_nclk_0.nRST PFD_0.VDD 0.60215f
C15 a_53065_20179# PFD_0.VDD 0.42601f
C16 a_64383_23434# 3bit_freq_divider_1.dff_nclk_0.D 0.0175f
C17 3bit_freq_divider_0.A0 m3_17285_2698# 0.30224f
C18 a_57178_43159# a_57084_43159# 0.42552f
C19 3bit_freq_divider_0.dff_nclk_0.nCLK a_53968_23946# 0.32517f
C20 a_54747_49259# charge_pump_0.vout 0.13589f
C21 a_45451_28860# PFD_0.VCO_CLK 0.12714f
C22 a_53022_43738# a_53058_43159# 0.24146f
C23 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.EN 0.12847f
C24 m2_16847_2260# m3_16847_2260# 0.2063p
C25 PFD_0.VDD a_53065_21935# 0.43552f
C26 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D PFD_0.VDD 0.97083f
C27 3bit_freq_divider_0.freq_div_cell_0.Cin 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.22232f
C28 a_60584_24580# a_60385_24717# 0.14868f
C29 3bit_freq_divider_1.freq_div_cell_0.Cin PFD_0.VDD 1.21632f
C30 a_53022_43738# a_53086_40850# 0.06371f
C31 a_61707_21488# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 0.24715f
C32 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.60301f
C33 3bit_freq_divider_1.sg13g2_or3_1_0.C a_63255_25000# 0.23357f
C34 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ 0.02712f
C35 a_57173_40413# a_58515_40413# 1.04202f
C36 a_58653_42591# a_58520_43159# 0.2448f
C37 a_54898_21129# a_54434_21392# 0.0104f
C38 a_54472_21129# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.12185f
C39 PFD_0.VDD a_53738_22270# 0.21577f
C40 a_61691_22290# a_61394_21976# 0.17766f
C41 a_53022_43738# a_57084_43159# 0.19696f
C42 a_61707_25000# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 0.24715f
C43 a_54842_49733# charge_pump_0.vout 0.02265f
C44 3bit_freq_divider_0.sg13g2_or3_1_0.C 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.05745f
C45 a_61707_25000# 3bit_freq_divider_1.freq_div_cell_0.Cin 0.01154f
C46 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_1.freq_div_cell_0.Cout 0.3426f
C47 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 0.40308f
C48 m6_16847_2260# m5_16847_2260# 0.13106p
C49 a_54472_24641# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.02559f
C50 a_61691_22290# PFD_0.VDD 0.68813f
C51 11Stage_vco_new_0.vctl a_54489_40413# 0.03623f
C52 a_56038_24617# a_56013_24979# 0.01952f
C53 a_51648_24041# a_51693_23075# 0.03957f
C54 a_51693_23075# a_51684_22692# 0.66077f
C55 a_64383_23889# a_64383_23628# 0.02302f
C56 3bit_freq_divider_1.A0 m5_17331_2744# 0.40842f
C57 a_62654_21971# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 0.01984f
C58 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.60301f
C59 3bit_freq_divider_0.sg13g2_nand2_1_0.Y PFD_0.VDD 3.38843f
C60 11Stage_vco_new_0.vctl a_55969_42591# 0.0811f
C61 11Stage_vco_new_0.vctl a_53152_43159# 0.01896f
C62 PFD_0.Ref_CLK a_45451_28860# 0.13923f
C63 a_51622_24863# PFD_0.VCO_CLK 0.02673f
C64 a_54489_40413# PFD_0.VDD 1.24454f
C65 a_62654_21971# 3bit_freq_divider_1.A2 0.02368f
C66 a_60967_23234# 3bit_freq_divider_1.freq_div_cell_0.Cout 0.13167f
C67 a_62270_24055# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.17312f
C68 a_64383_23706# PFD_0.VDD 0.30655f
C69 3bit_freq_divider_0.dff_nclk_0.nRST 3bit_freq_divider_0.A0 0.14477f
C70 a_54494_43159# a_55742_43159# 0.10125f
C71 3bit_freq_divider_0.freq_div_cell_0.Cin a_54472_22885# 0.01011f
C72 a_55969_42591# PFD_0.VDD 0.0108f
C73 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_0.Cin 0.32366f
C74 a_53152_43159# PFD_0.VDD 1.21324f
C75 a_64384_21091# a_64714_21414# 0.014f
C76 a_61887_22290# a_62119_22361# 0.13068f
C77 a_64383_23706# 3bit_freq_divider_1.dff_nclk_0.D 0.12409f
C78 a_58453_40283# a_57173_40413# 0.45932f
C79 3bit_freq_divider_0.CLK_IN 3bit_freq_divider_0.EN 0.41907f
C80 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 3bit_freq_divider_1.dff_nclk_0.nCLK 0.02503f
C81 a_62900_23691# 3bit_freq_divider_1.A2 0.01917f
C82 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_51684_22692# 0.01473f
C83 a_64383_23434# a_64419_23326# 0.66077f
C84 3bit_freq_divider_0.dff_nclk_0.D a_51684_22284# 0.43097f
C85 3bit_freq_divider_0.dff_nclk_0.D PFD_0.VCO_CLK 0.01884f
C86 a_62654_21971# PFD_0.VDD 0.4336f
C87 a_60385_24717# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI 0.02161f
C88 3bit_freq_divider_0.sg13g2_or3_1_0.C a_51648_21103# 0.25034f
C89 a_54427_40283# a_54489_40413# 0.12319f
C90 a_53774_20178# a_53968_20434# 0.05314f
C91 a_53065_20179# a_53899_20488# 0.03957f
C92 a_53738_24026# a_53968_23946# 0.13068f
C93 a_61707_21488# 3bit_freq_divider_1.freq_div_cell_0.Cout 0.12082f
C94 3bit_freq_divider_1.freq_div_cell_0.Cout 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 0.084f
C95 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.sg13g2_or3_1_0.C 0.13894f
C96 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_0.freq_div_cell_0.Cin 0.084f
C97 3bit_freq_divider_1.CLK_OUT m7_16847_2260# 1.40976f
C98 3bit_freq_divider_1.dff_nclk_0.nRST 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.16234f
C99 a_62900_23691# PFD_0.VDD 0.31029f
C100 11Stage_vco_new_0.vctl 3bit_freq_divider_0.CLK_IN 0.4797f
C101 a_63255_23244# a_63426_22886# 0.36535f
C102 a_64383_23300# PFD_0.VDD 0.29403f
C103 a_64424_22200# 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.0838f
C104 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.A2 0.64366f
C105 3bit_freq_divider_1.A2 a_63255_21488# 0.39947f
C106 a_46749_30782# a_47777_29803# 0.4544f
C107 3bit_freq_divider_0.dff_nclk_0.nCLK a_53899_22244# 0.17328f
C108 3bit_freq_divider_1.A1 3bit_freq_divider_1.CLK_OUT 0.01478f
C109 3bit_freq_divider_0.CLK_IN PFD_0.VDD 2.00225f
C110 a_64383_23300# 3bit_freq_divider_1.dff_nclk_0.D 0.04146f
C111 a_61394_23732# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 0.3562f
C112 a_57173_40413# a_57112_40850# 0.03198f
C113 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.21745f
C114 a_53022_43738# a_57173_40413# 0.05042f
C115 3bit_freq_divider_0.dff_nclk_0.nCLK a_52924_22885# 0.03415f
C116 a_54898_24641# a_54434_24904# 0.0104f
C117 a_54472_24641# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 0.12185f
C118 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ a_53445_20214# 0.10118f
C119 3bit_freq_divider_1.A0 a_63255_25000# 0.39999f
C120 a_54504_22015# a_53738_22270# 0.47248f
C121 a_51693_23075# a_51631_22774# 0.04255f
C122 PFD_0.VDD a_63255_21488# 0.26051f
C123 a_51622_24863# a_51721_24988# 0.0229f
C124 a_61707_21488# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 0.46099f
C125 a_61691_22290# a_62119_22361# 0.05314f
C126 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.dff_nclk_0.D 0.04354f
C127 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_1.A2 0.20327f
C128 a_56013_24979# a_56137_24678# 0.10864f
C129 a_52886_23148# 3bit_freq_divider_0.A1 0.39847f
C130 sg13g2_inv_1_0.A 3bit_freq_divider_0.EN 0.24728f
C131 a_52950_23913# PFD_0.VDD 0.24052f
C132 3bit_freq_divider_1.sg13g2_nand2_1_0.Y a_60967_23234# 0.08797f
C133 a_51693_23075# 3bit_freq_divider_0.A1 0.01284f
C134 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI 0.42892f
C135 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_52924_24641# 0.02246f
C136 a_51693_23075# a_51693_23426# 0.70262f
C137 3bit_freq_divider_1.A1 a_63426_24642# 0.01474f
C138 a_53152_43159# a_53285_42591# 0.22422f
C139 PFD_0.VCO_CLK a_46817_27899# 0.92547f
C140 3bit_freq_divider_0.sg13g2_nand2_1_0.Y a_55345_21385# 0.08797f
C141 a_48909_28913# a_47954_28913# 0.39061f
C142 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.60301f
C143 3bit_freq_divider_0.EN PFD_0.VDD 6.40652f
C144 PFD_0.VDD a_53774_21934# 0.69275f
C145 a_55836_43159# a_57178_43159# 1.16874f
C146 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ PFD_0.VDD 0.18065f
C147 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q PFD_0.VDD 1.41895f
C148 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_52886_24904# 0.14987f
C149 3bit_freq_divider_1.CLK_OUT m4_17285_2698# 0.3817f
C150 a_51685_23725# 3bit_freq_divider_0.dff_nclk_0.D 0.12409f
C151 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_51631_22774# 0.33833f
C152 a_53022_43738# a_57111_40283# 0.18962f
C153 m3_16847_2260# m4_16847_2260# 0.2063p
C154 PFD_0.VDD 3bit_freq_divider_1.A2 1.18034f
C155 a_51648_21103# a_51708_21299# 0.02055f
C156 a_62119_24117# PFD_0.VDD 0.32287f
C157 3bit_freq_divider_1.A2 3bit_freq_divider_1.sg13g2_or3_1_0.B 0.1586f
C158 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 0.05125f
C159 a_51759_25014# PFD_0.VDD 0.0834f
C160 a_63426_21130# a_63255_21488# 0.36535f
C161 11Stage_vco_new_0.vctl PFD_0.VDD 0.29003f
C162 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_0.A1 0.15458f
C163 a_62654_20215# a_63463_20216# 0.09575f
C164 3bit_freq_divider_0.A1 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.02018f
C165 sg13g2_inv_1_0.A PFD_0.VDD 3.87548f
C166 a_54434_24904# PFD_0.VDD 0.27564f
C167 a_61394_21976# PFD_0.VDD 0.38024f
C168 a_54400_43159# a_53152_43159# 0.09095f
C169 a_53022_43738# a_55836_43159# 0.05231f
C170 a_51648_24041# 3bit_freq_divider_0.dff_nclk_0.nRST 0.30513f
C171 a_51684_22692# 3bit_freq_divider_0.dff_nclk_0.nRST 0.126f
C172 a_61691_24046# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.35198f
C173 a_53445_20214# a_53738_20514# 0.04306f
C174 a_64383_23300# a_64419_23326# 0.70262f
C175 3bit_freq_divider_1.freq_div_cell_1.Cout 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 0.04623f
C176 3bit_freq_divider_0.EN charge_pump_0.bias_n 0.02661f
C177 a_57178_43159# a_58653_42591# 0.03197f
C178 3bit_freq_divider_1.A1 m5_17331_2744# 0.40842f
C179 PFD_0.VDD 3bit_freq_divider_1.sg13g2_or3_1_0.B 0.10974f
C180 a_64362_24865# a_64398_24796# 0.14868f
C181 3bit_freq_divider_1.A1 3bit_freq_divider_1.dff_nclk_0.nCLK 0.23798f
C182 a_52944_43077# a_53147_40413# 0.83377f
C183 PFD_0.VDD 3bit_freq_divider_1.dff_nclk_0.D 0.84615f
C184 3bit_freq_divider_1.dff_nclk_0.nRST a_64362_24865# 0.03098f
C185 a_51648_24438# PFD_0.VCO_CLK 0.11636f
C186 a_62654_23727# a_62900_23691# 0.41048f
C187 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 0.22983f
C188 a_54434_23148# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 0.24715f
C189 3bit_freq_divider_0.EN 3bit_freq_divider_0.A0 0.11772f
C190 a_61707_25000# PFD_0.VDD 0.27566f
C191 a_63426_21130# 3bit_freq_divider_1.A2 0.02209f
C192 a_54427_40283# PFD_0.VDD 1.36601f
C193 PFD_0.VDD a_52924_21129# 0.20953f
C194 a_55948_56737# charge_pump_0.bias_p 0.02673f
C195 sg13g2_inv_1_0.A charge_pump_0.bias_n 0.06869f
C196 3bit_freq_divider_1.sg13g2_or3_1_0.C 3bit_freq_divider_1.A0 0.12518f
C197 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.40308f
C198 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_53065_20179# 0.01984f
C199 PFD_0.VDD charge_pump_0.bias_n 0.83592f
C200 a_53445_23726# PFD_0.VDD 0.31261f
C201 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_53065_21935# 0.0119f
C202 a_63426_21130# PFD_0.VDD 0.20953f
C203 3bit_freq_divider_0.dff_nclk_0.nCLK a_53968_20434# 0.32507f
C204 a_62270_20543# a_62654_20215# 0.03957f
C205 a_47954_28913# PFD_0.VDD 0.45155f
C206 PFD_0.VDD a_61691_20534# 0.67211f
C207 a_58520_43159# 3bit_freq_divider_0.CLK_IN 0.83486f
C208 m5_17331_2744# m4_17285_2698# 0.1814p
C209 11Stage_vco_new_0.vctl a_59800_40852# 0.05123f
C210 PFD_0.Ref_CLK m7_16847_2260# 1.44946f
C211 a_58734_56203# a_58536_54976# 0.19076f
C212 PFD_0.DOWN PFD_0.VDD 1.56226f
C213 a_53774_21934# a_54504_22015# 0.17766f
C214 11Stage_vco_new_0.vctl a_53285_42591# 0.08086f
C215 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VDD 0.27798f
C216 3bit_freq_divider_1.CLK_OUT a_64398_24796# 0.02652f
C217 3bit_freq_divider_0.freq_div_cell_1.Cout 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.04623f
C218 PFD_0.VDD 3bit_freq_divider_0.A0 1.32697f
C219 a_64383_23434# 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01473f
C220 a_54504_20259# PFD_0.VDD 0.36995f
C221 3bit_freq_divider_1.dff_nclk_0.nRST 3bit_freq_divider_1.CLK_OUT 0.07748f
C222 3bit_freq_divider_1.freq_div_cell_1.Cout 3bit_freq_divider_1.freq_div_cell_0.Cout 0.09134f
C223 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 0.22983f
C224 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_0.Cin 0.22232f
C225 a_62654_23727# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 0.0119f
C226 3bit_freq_divider_0.sg13g2_or3_1_0.B PFD_0.VDD 0.11082f
C227 3bit_freq_divider_0.dff_nclk_0.nRST a_51631_22774# 0.3267f
C228 3bit_freq_divider_1.A1 a_63255_25000# 0.01849f
C229 a_61394_21976# a_62119_22361# 0.45825f
C230 a_61394_23732# a_62119_24117# 0.45825f
C231 a_53899_20488# PFD_0.VDD 0.24492f
C232 a_53774_23690# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.33731f
C233 PFD_0.VDD a_64419_23326# 0.2446f
C234 a_62900_23691# a_61887_24046# 0.04306f
C235 a_62654_23727# 3bit_freq_divider_1.A2 0.02178f
C236 a_60385_24947# a_60584_24580# 0.0229f
C237 3bit_freq_divider_1.dff_nclk_0.nCLK a_63463_20216# 0.05882f
C238 a_53085_40283# a_53147_40413# 0.104f
C239 a_57173_40413# a_55831_40413# 1.08982f
C240 a_62119_22361# PFD_0.VDD 0.31854f
C241 3bit_freq_divider_0.A1 3bit_freq_divider_0.dff_nclk_0.nRST 0.08188f
C242 3bit_freq_divider_0.sg13g2_or3_1_0.C 3bit_freq_divider_0.A2 0.04643f
C243 a_51693_23426# 3bit_freq_divider_0.dff_nclk_0.nRST 0.3148f
C244 a_53774_20178# a_53738_20514# 0.44698f
C245 PFD_0.VDD a_55345_21385# 0.45855f
C246 3bit_freq_divider_1.dff_nclk_0.D a_64419_23326# 0.01591f
C247 a_54434_23148# 3bit_freq_divider_0.freq_div_cell_0.Cout 0.01154f
C248 PFD_0.VDD a_54504_22015# 0.38024f
C249 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_0.Cout 0.22232f
C250 PFD_0.DOWN charge_pump_0.bias_n 0.01578f
C251 3bit_freq_divider_1.freq_div_cell_0.Cout a_61707_23244# 0.01154f
C252 a_61394_23732# PFD_0.VDD 0.38531f
C253 a_63463_23728# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 0.21609f
C254 a_61887_20534# a_62119_20605# 0.13068f
C255 11Stage_vco_new_0.vctl a_58520_43159# 0.20162f
C256 a_62654_23727# PFD_0.VDD 0.43765f
C257 a_61887_20534# a_62270_20543# 0.66077f
C258 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_20534# 0.33731f
C259 3bit_freq_divider_1.A1 a_63426_22886# 0.01971f
C260 3bit_freq_divider_1.freq_div_cell_1.Cout 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 0.2223f
C261 a_61878_22886# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 0.12185f
C262 a_55345_24897# PFD_0.VDD 0.45478f
C263 a_54400_43159# PFD_0.VDD 1.37065f
C264 a_64384_21091# a_64714_21300# 0.02055f
C265 PFD_0.Ref_CLK m4_17285_2698# 0.39515f
C266 PFD_0.Ref_CLK a_47777_29803# 0.17902f
C267 a_45579_29803# a_46749_30782# 0.25388f
C268 a_64459_24995# a_64362_24865# 0.10864f
C269 sg13g2_inv_1_0.A a_56742_53480# 0.28042f
C270 a_60967_21478# 3bit_freq_divider_1.freq_div_cell_0.Cout 0.13034f
C271 a_58520_43159# PFD_0.VDD 1.48446f
C272 a_54434_24904# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 0.12082f
C273 a_61707_25000# a_61675_24642# 0.0104f
C274 a_54504_23771# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.08213f
C275 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.1064f
C276 a_53065_20179# a_53445_20214# 0.41048f
C277 a_64384_21091# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.33258f
C278 a_58426_43159# PFD_0.VDD 1.37111f
C279 a_57111_40283# a_55831_40413# 0.45742f
C280 PFD_0.VDD 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 0.77158f
C281 a_58515_40413# 3bit_freq_divider_0.CLK_IN 0.04768f
C282 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_0.CLK_IN 0.02001f
C283 3bit_freq_divider_1.dff_nclk_0.nCLK a_62119_20605# 0.32732f
C284 a_64384_24445# PFD_0.VDD 0.24105f
C285 3bit_freq_divider_1.freq_div_cell_1.Cout 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.07626f
C286 3bit_freq_divider_1.dff_nclk_0.nCLK a_62270_20543# 0.17248f
C287 a_52886_21392# PFD_0.VDD 0.26051f
C288 a_56013_24979# PFD_0.VDD 0.11379f
C289 a_61887_24046# a_62119_24117# 0.13068f
C290 a_51648_21103# 3bit_freq_divider_0.sg13g2_or3_1_0.A 0.31317f
C291 a_64384_24445# 3bit_freq_divider_1.dff_nclk_0.D 0.2233f
C292 a_52944_43077# a_53085_40283# 0.45412f
C293 3bit_freq_divider_1.dff_nclk_0.nRST a_64383_23628# 0.3268f
C294 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ a_62900_20179# 0.10118f
C295 PFD_0.Ref_CLK m1_17285_2698# 0.01061f
C296 PFD_0.VDD a_54434_21392# 0.2676f
C297 a_54494_43159# a_55836_43159# 1.11028f
C298 a_64383_23628# a_64424_22200# 0.17766f
C299 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.sg13g2_or3_1_0.A 0.48568f
C300 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_60967_21478# 0.30546f
C301 a_56742_53480# charge_pump_0.bias_n 0.05592f
C302 a_59097_54704# charge_pump_0.bias_p 0.04726f
C303 3bit_freq_divider_1.CLK_OUT m3_17285_2698# 0.2919f
C304 a_55345_23141# 3bit_freq_divider_0.freq_div_cell_0.Cout 0.13167f
C305 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 0.05125f
C306 a_53899_24000# a_53774_23690# 0.04304f
C307 3bit_freq_divider_1.A1 3bit_freq_divider_1.sg13g2_or3_1_0.C 0.16352f
C308 a_61887_24046# PFD_0.VDD 0.22153f
C309 a_55941_24882# a_56137_24678# 0.0229f
C310 a_52886_21392# a_52924_21129# 0.36535f
C311 a_51648_24041# PFD_0.VDD 0.41893f
C312 3bit_freq_divider_0.sg13g2_or3_1_0.C a_52924_24641# 0.10662f
C313 a_53022_43738# a_54489_40413# 0.06435f
C314 a_51684_22692# PFD_0.VDD 0.19308f
C315 a_55831_40413# a_55770_40850# 0.03239f
C316 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ 0.08555f
C317 a_54357_49278# PFD_0.VDD 0.31963f
C318 a_60385_24717# PFD_0.VDD 0.11381f
C319 a_55862_56737# PFD_0.VDD 0.47223f
C320 a_53086_40850# a_53147_40413# 0.0531f
C321 a_61887_22290# a_62270_22299# 0.66077f
C322 a_62900_21935# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.27425f
C323 a_58520_43159# a_59800_40852# 0.12912f
C324 a_53022_43738# a_53152_43159# 0.08528f
C325 PFD_0.VDD a_62900_20179# 0.30479f
C326 3bit_freq_divider_1.freq_div_cell_1.Cout a_61707_21488# 0.01154f
C327 a_55836_43159# a_57311_42591# 0.03197f
C328 3bit_freq_divider_0.sg13g2_or3_1_0.C a_52886_24904# 0.23357f
C329 3bit_freq_divider_1.sg13g2_nand2_1_0.Y a_60967_21478# 0.08797f
C330 11Stage_vco_new_0.vctl a_58515_40413# 0.02252f
C331 3bit_freq_divider_0.dff_nclk_0.nCLK a_53968_22190# 0.32534f
C332 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q PFD_0.VDD 1.42261f
C333 3bit_freq_divider_1.A1 a_63463_23728# 0.03561f
C334 a_58515_40413# PFD_0.VDD 1.43082f
C335 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_63463_20216# 0.12389f
C336 a_51684_22284# 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.0838f
C337 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_1.A2 0.21293f
C338 3bit_freq_divider_1.A1 a_63255_23244# 0.39563f
C339 a_55862_56737# charge_pump_0.bias_n 0.34812f
C340 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.1064f
C341 a_61707_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 0.24715f
C342 a_53065_20179# a_53774_20178# 0.02335f
C343 a_52950_20401# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ 0.21609f
C344 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.sg13g2_or3_1_0.A 0.48568f
C345 3bit_freq_divider_0.A1 3bit_freq_divider_0.EN 0.5347f
C346 a_51648_24041# 3bit_freq_divider_0.A0 0.0271f
C347 a_54357_49278# PFD_0.DOWN 0.04759f
C348 3bit_freq_divider_0.dff_nclk_0.nCLK a_52886_23148# 0.10223f
C349 PFD_0.UP PFD_0.VDD 0.82664f
C350 3bit_freq_divider_0.dff_nclk_0.nCLK a_53738_20514# 0.18358f
C351 a_61691_20534# a_62900_20179# 0.04324f
C352 a_45658_27900# PFD_0.VDD 1.00659f
C353 a_59600_42432# 3bit_freq_divider_0.CLK_IN 0.01283f
C354 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q PFD_0.VDD 1.66358f
C355 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_52924_21129# 0.01011f
C356 a_61691_22290# a_62270_22299# 0.04304f
C357 a_53058_43159# a_52944_43077# 0.09058f
C358 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_0.Cout 0.3426f
C359 a_55345_24897# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 0.21784f
C360 11Stage_vco_new_0.vctl charge_pump_0.vout 0.05724f
C361 a_52944_43077# a_53086_40850# 0.23665f
C362 PFD_0.VDD 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.28742f
C363 a_58426_43159# a_58520_43159# 0.4131f
C364 a_53065_23691# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 0.0119f
C365 3bit_freq_divider_1.A0 m7_16847_2260# 1.40976f
C366 PFD_0.VDD a_51631_22774# 0.62631f
C367 a_61878_24642# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI 0.01011f
C368 a_53065_23691# a_53774_23690# 0.02335f
C369 a_52950_23913# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ 0.21609f
C370 a_58453_40283# PFD_0.VDD 1.38336f
C371 3bit_freq_divider_1.dff_nclk_0.D 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.17618f
C372 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_61707_25000# 0.46099f
C373 charge_pump_0.vout PFD_0.VDD 0.06128f
C374 11Stage_vco_new_0.vctl a_57178_43159# 0.02155f
C375 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_54472_22885# 0.02559f
C376 a_54434_23148# a_54472_22885# 0.36535f
C377 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 1.03924f
C378 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D a_53774_21934# 0.01446f
C379 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.10701f
C380 3bit_freq_divider_0.A1 PFD_0.VDD 1.47452f
C381 a_61394_23732# a_61887_24046# 0.47248f
C382 3bit_freq_divider_1.A1 3bit_freq_divider_1.A0 1.97044f
C383 a_61691_24046# a_62270_24055# 0.04304f
C384 a_51693_23426# PFD_0.VDD 0.29403f
C385 3bit_freq_divider_0.dff_nclk_0.nCLK a_53774_23690# 0.35198f
C386 a_62654_23727# a_61887_24046# 0.40027f
C387 a_57178_43159# PFD_0.VDD 1.6124f
C388 3bit_freq_divider_0.dff_nclk_0.D a_51648_24438# 0.2233f
C389 a_62270_22299# a_62654_21971# 0.03957f
C390 3bit_freq_divider_0.EN a_58536_54976# 0.21462f
C391 a_58515_40413# a_59800_40852# 0.21632f
C392 a_61887_22290# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.18493f
C393 a_56013_24979# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 0.02161f
C394 11Stage_vco_new_0.vctl a_57112_40850# 0.05026f
C395 3bit_freq_divider_1.dff_nclk_0.nRST a_64731_24890# 0.01267f
C396 a_53022_43738# 11Stage_vco_new_0.vctl 0.09064f
C397 PFD_0.DOWN PFD_0.UP 0.20773f
C398 a_52924_24641# a_52886_24904# 0.36535f
C399 PFD_0.DOWN a_45658_27900# 0.61911f
C400 3bit_freq_divider_0.dff_nclk_0.nCLK a_53445_21970# 0.27428f
C401 3bit_freq_divider_1.A1 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 0.01108f
C402 a_61394_20220# a_62119_20605# 0.45825f
C403 a_60385_24558# PFD_0.VDD 0.04481f
C404 3bit_freq_divider_1.sg13g2_or3_1_0.C a_64384_21091# 0.25034f
C405 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D a_53774_23690# 0.01446f
C406 charge_pump_0.vout charge_pump_0.bias_n 0.23558f
C407 a_61878_22886# a_61707_23244# 0.36535f
C408 a_53022_43738# PFD_0.VDD 13.1748f
C409 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 0.97883f
C410 a_62900_21935# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ 0.10118f
C411 PFD_0.Ref_CLK m3_17285_2698# 0.30224f
C412 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_55345_21385# 0.30546f
C413 a_64383_23434# a_64383_23628# 0.44985f
C414 PFD_0.Ref_CLK a_45579_29803# 1.21724f
C415 a_53445_20214# PFD_0.VDD 0.30479f
C416 3bit_freq_divider_1.dff_nclk_0.nRST 3bit_freq_divider_1.sg13g2_or3_1_0.C 0.57774f
C417 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ PFD_0.VDD 0.18755f
C418 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_1.dff_nclk_0.nCLK 0.21603f
C419 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.dff_nclk_0.nCLK 0.32366f
C420 a_51684_22284# 3bit_freq_divider_0.dff_nclk_0.nRST 0.34874f
C421 3bit_freq_divider_1.A0 m4_17285_2698# 0.3817f
C422 PFD_0.VCO_CLK 3bit_freq_divider_0.dff_nclk_0.nRST 0.06912f
C423 PFD_0.VDD a_58536_54976# 0.98046f
C424 3bit_freq_divider_0.dff_nclk_0.nCLK a_54504_23771# 0.37259f
C425 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ 0.08742f
C426 a_61887_22290# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01324f
C427 a_53022_43738# a_54427_40283# 0.19046f
C428 a_55769_40283# a_54489_40413# 0.45471f
C429 3bit_freq_divider_0.A1 3bit_freq_divider_0.A0 0.55463f
C430 a_54489_40413# a_55831_40413# 1.05293f
C431 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_53738_20514# 0.01324f
C432 a_58515_40413# a_58520_43159# 1.39948f
C433 a_61691_22290# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.35569f
C434 3bit_freq_divider_0.A2 3bit_freq_divider_0.sg13g2_or3_1_0.A 0.2051f
C435 m6_17427_2840# 3bit_freq_divider_0.A0 1.23795f
C436 3bit_freq_divider_0.A1 3bit_freq_divider_0.sg13g2_or3_1_0.B 0.27832f
C437 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_62654_23727# 0.02071f
C438 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D a_54504_23771# 0.3562f
C439 a_51648_24041# a_51684_22692# 0.40027f
C440 a_46749_30782# PFD_0.VDD 1.12191f
C441 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ a_62654_20215# 0.0571f
C442 a_54494_43159# a_55969_42591# 0.03197f
C443 a_53738_24026# a_53774_23690# 0.44698f
C444 a_53445_23726# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ 0.10118f
C445 a_64362_24865# PFD_0.VDD 0.08341f
C446 a_53152_43159# a_54494_43159# 1.07553f
C447 a_61691_24046# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.33731f
C448 3bit_freq_divider_0.dff_nclk_0.nCLK a_52950_22157# 0.05957f
C449 a_58536_54976# charge_pump_0.bias_n 0.02549f
C450 a_58734_56203# charge_pump_0.bias_p 0.03822f
C451 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VDD 0.30706f
C452 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_52886_21392# 0.12248f
C453 a_53968_23946# a_53774_23690# 0.05314f
C454 a_54489_40413# a_54428_40850# 0.03832f
C455 a_53022_43738# a_59800_40852# 0.01439f
C456 3bit_freq_divider_0.dff_nclk_0.nCLK a_53065_20179# 0.31132f
C457 a_64383_23628# a_64383_23706# 0.04324f
C458 a_55941_24882# PFD_0.VDD 0.10494f
C459 a_61878_24642# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 0.12185f
C460 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_54434_21392# 0.46099f
C461 a_62654_21971# a_63463_21972# 0.09575f
C462 a_62654_21971# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.31887f
C463 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_0.Cout 1.22849f
C464 a_53022_43738# a_53285_42591# 0.02036f
C465 a_61691_22290# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.33731f
C466 3bit_freq_divider_0.dff_nclk_0.nCLK a_53065_21935# 0.31904f
C467 PFD_0.VDD a_62654_20215# 0.42601f
C468 a_62270_22299# PFD_0.VDD 0.26052f
C469 a_53899_22244# a_53968_22190# 0.70262f
C470 a_64383_23889# 3bit_freq_divider_1.dff_nclk_0.nRST 0.30513f
C471 a_62900_23691# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.24211f
C472 3bit_freq_divider_1.A1 m7_16847_2260# 1.40976f
C473 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D a_54504_22015# 0.3562f
C474 3bit_freq_divider_0.dff_nclk_0.nCLK a_53738_22270# 0.18642f
C475 a_53738_24026# a_54504_23771# 0.47248f
C476 a_57178_43159# a_58520_43159# 0.20611f
C477 a_51685_23725# 3bit_freq_divider_0.dff_nclk_0.nRST 0.25925f
C478 a_63223_24642# a_63255_25000# 0.0104f
C479 m1_17285_2698# m2_17285_2698# 0.20496p
C480 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.freq_div_cell_0.Cout 0.10559f
C481 3bit_freq_divider_0.sg13g2_or3_1_0.C a_51693_23075# 0.01089f
C482 3bit_freq_divider_1.CLK_OUT PFD_0.VDD 0.38178f
C483 a_53774_20178# PFD_0.VDD 0.67672f
C484 a_53968_23946# a_54504_23771# 0.45825f
C485 a_57178_43159# a_58426_43159# 0.09524f
C486 3bit_freq_divider_1.freq_div_cell_1.Cout a_60967_21478# 0.13166f
C487 a_54357_49278# PFD_0.UP 0.30851f
C488 a_48909_28913# PFD_0.VCO_CLK 0.1514f
C489 a_64383_23300# a_64383_23628# 0.05314f
C490 3bit_freq_divider_0.freq_div_cell_0.Cin 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 0.42266f
C491 3bit_freq_divider_0.freq_div_cell_0.Cin a_54434_23148# 0.12082f
C492 a_53022_43738# a_54400_43159# 0.19723f
C493 3bit_freq_divider_1.CLK_OUT 3bit_freq_divider_1.dff_nclk_0.D 0.01884f
C494 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.23907f
C495 a_52950_20401# a_53065_20179# 0.09575f
C496 a_53022_43738# a_58520_43159# 0.15068f
C497 3bit_freq_divider_1.dff_nclk_0.nCLK a_63255_21488# 0.10313f
C498 a_61878_21130# PFD_0.VDD 0.21321f
C499 a_52886_23148# a_52924_22885# 0.36535f
C500 a_61691_20534# a_62654_20215# 0.02302f
C501 a_59600_42432# a_58520_43159# 0.01604f
C502 a_51648_24041# a_51631_22774# 0.02302f
C503 a_51684_22692# a_51631_22774# 0.45006f
C504 a_60385_24947# PFD_0.VDD 0.11858f
C505 a_63426_24642# PFD_0.VDD 0.20944f
C506 a_53022_43738# a_58426_43159# 0.10045f
C507 3bit_freq_divider_0.sg13g2_or3_1_0.C 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.28129f
C508 a_54357_49278# charge_pump_0.vout 0.01432f
C509 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.04726f
C510 PFD_0.VDD a_61887_20534# 0.19386f
C511 11Stage_vco_new_0.vctl a_55831_40413# 0.03134f
C512 3bit_freq_divider_0.A1 a_51684_22692# 0.03873f
C513 3bit_freq_divider_0.dff_nclk_0.D a_51693_23075# 0.01591f
C514 a_51693_23426# a_51684_22692# 0.13068f
C515 a_53899_24000# PFD_0.VDD 0.26493f
C516 a_63463_21972# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 0.12389f
C517 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ 3bit_freq_divider_1.dff_nclk_0.nCLK 0.08552f
C518 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_1.dff_nclk_0.nCLK 1.03922f
C519 a_52950_23913# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.12519f
C520 a_55769_40283# PFD_0.VDD 1.36975f
C521 11Stage_vco_new_0.vctl a_54494_43159# 0.02166f
C522 PFD_0.Ref_CLK a_48909_28913# 0.12375f
C523 a_45579_29803# a_45451_28860# 0.44406f
C524 a_55831_40413# PFD_0.VDD 1.18769f
C525 a_64383_23434# 3bit_freq_divider_1.sg13g2_or3_1_0.C 0.03556f
C526 a_63463_21972# 3bit_freq_divider_1.A2 0.01788f
C527 3bit_freq_divider_1.A1 m4_17285_2698# 0.3817f
C528 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.A2 0.86741f
C529 a_62119_24117# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.32742f
C530 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_52924_22885# 0.01011f
C531 a_64714_21300# PFD_0.VDD 0.01263f
C532 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 3bit_freq_divider_0.EN 0.02092f
C533 a_54472_21129# PFD_0.VDD 0.21321f
C534 a_55836_43159# a_55742_43159# 0.42065f
C535 a_55345_21385# 3bit_freq_divider_0.freq_div_cell_0.Cout 0.13034f
C536 a_54504_20259# a_53774_20178# 0.17766f
C537 a_54494_43159# PFD_0.VDD 1.48562f
C538 a_62270_22299# a_62119_22361# 0.70262f
C539 a_61394_21976# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.37259f
C540 a_58453_40283# a_58515_40413# 0.1135f
C541 a_60385_24558# a_60385_24717# 0.01952f
C542 11Stage_vco_new_0.vctl a_54428_40850# 0.04894f
C543 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.04726f
C544 3bit_freq_divider_0.dff_nclk_0.D 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.17618f
C545 a_63463_21972# PFD_0.VDD 0.2345f
C546 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.25573f
C547 PFD_0.VDD 3bit_freq_divider_1.dff_nclk_0.nCLK 2.89514f
C548 a_53774_20178# a_53899_20488# 0.04304f
C549 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.sg13g2_or3_1_0.B 0.58488f
C550 a_52950_23913# a_53065_23691# 0.09575f
C551 3bit_freq_divider_0.freq_div_cell_0.Cin a_55345_23141# 0.13034f
C552 11Stage_vco_new_0.vctl a_57311_42591# 0.08436f
C553 a_54434_24904# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.46099f
C554 a_61691_20534# a_61887_20534# 0.45047f
C555 3bit_freq_divider_1.dff_nclk_0.D 3bit_freq_divider_1.dff_nclk_0.nCLK 0.04354f
C556 PFD_0.VDD a_54428_40850# 0.01482f
C557 a_62654_21971# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ 0.0571f
C558 a_64383_23628# PFD_0.VDD 0.62587f
C559 a_51684_22284# PFD_0.VDD 0.36995f
C560 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61887_20534# 0.01324f
C561 PFD_0.VCO_CLK PFD_0.VDD 1.82327f
C562 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q PFD_0.VDD 1.68952f
C563 3bit_freq_divider_1.freq_div_cell_0.Cin a_60967_23234# 0.13034f
C564 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D PFD_0.VDD 0.9437f
C565 PFD_0.Ref_CLK 3bit_freq_divider_0.EN 0.09396f
C566 a_64383_23628# 3bit_freq_divider_1.dff_nclk_0.D 0.03728f
C567 m4_16847_2260# m5_16847_2260# 0.2063p
C568 a_62654_21971# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 0.0119f
C569 a_55941_24882# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 0.12404f
C570 a_56695_49467# charge_pump_0.vout 0.02916f
C571 3bit_freq_divider_1.A0 m3_17285_2698# 0.2919f
C572 a_61394_21976# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.08213f
C573 3bit_freq_divider_0.dff_nclk_0.nCLK a_53774_21934# 0.35569f
C574 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.10521f
C575 a_57173_40413# a_58454_40850# 0.22936f
C576 a_53022_43738# a_58515_40413# 0.0744f
C577 a_56013_24979# a_55941_24882# 0.14868f
C578 a_53147_40413# a_54489_40413# 0.29213f
C579 3bit_freq_divider_0.A1 a_51631_22774# 0.02271f
C580 PFD_0.VDD 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.29872f
C581 a_63426_21130# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.03449f
C582 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_53738_22270# 0.01324f
C583 a_51693_23426# a_51631_22774# 0.05331f
C584 3bit_freq_divider_1.dff_nclk_0.nCLK a_61691_20534# 0.35517f
C585 a_63255_25000# 3bit_freq_divider_1.A2 0.02709f
C586 a_54434_21392# 3bit_freq_divider_0.freq_div_cell_0.Cout 0.12082f
C587 a_53065_23691# PFD_0.VDD 0.44373f
C588 m5_17331_2744# 3bit_freq_divider_0.A0 0.42278f
C589 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_0.Cout 0.22232f
C590 a_51648_21103# PFD_0.VDD 0.34051f
C591 3bit_freq_divider_0.sg13g2_or3_1_0.C 3bit_freq_divider_0.dff_nclk_0.nRST 0.57774f
C592 a_51693_23426# 3bit_freq_divider_0.A1 0.01735f
C593 3bit_freq_divider_0.CLK_IN 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 0.02001f
C594 a_64383_23434# a_64383_23889# 0.40027f
C595 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.dff_nclk_0.nCLK 0.60301f
C596 PFD_0.Ref_CLK PFD_0.VDD 2.49441f
C597 a_53738_20514# a_53968_20434# 0.13068f
C598 a_53152_43159# a_54627_42591# 0.03153f
C599 a_61878_24642# PFD_0.VDD 0.21401f
C600 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_1.Cout 0.07626f
C601 PFD_0.VCO_CLK a_47954_28913# 1.24436f
C602 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.11142f
C603 a_64384_24445# 3bit_freq_divider_1.CLK_OUT 0.1244f
C604 PFD_0.VDD a_54472_22885# 0.21321f
C605 3bit_freq_divider_0.dff_nclk_0.nCLK PFD_0.VDD 2.90191f
C606 m2_17285_2698# m3_17285_2698# 0.20496p
C607 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D a_61691_20534# 0.01446f
C608 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_63426_22886# 0.01011f
C609 a_63255_21488# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 0.12248f
C610 a_51759_25014# a_51721_24988# 0.10864f
C611 a_63255_25000# PFD_0.VDD 0.26507f
C612 a_61691_22290# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 0.01446f
C613 PFD_0.DOWN PFD_0.VCO_CLK 0.20401f
C614 a_51622_24863# 3bit_freq_divider_0.dff_nclk_0.nRST 0.10221f
C615 PFD_0.VCO_CLK 3bit_freq_divider_0.A0 0.1115f
C616 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_0.A0 0.24362f
C617 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.40308f
C618 3bit_freq_divider_0.freq_div_cell_0.Cin 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.25573f
C619 a_53022_43738# a_58453_40283# 0.19288f
C620 a_61878_24642# a_61707_25000# 0.36535f
C621 a_54434_24904# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 0.24715f
C622 a_53065_21935# a_53899_22244# 0.03957f
C623 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ 0.02712f
C624 a_51721_24988# PFD_0.VDD 0.08543f
C625 a_62119_22361# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.32758f
C626 PFD_0.VDD 3bit_freq_divider_1.freq_div_cell_0.Cout 1.22849f
C627 a_62654_20215# a_62900_20179# 0.41048f
C628 m6_16847_2260# m7_16847_2260# 39.787f
C629 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D PFD_0.VDD 0.97078f
C630 3bit_freq_divider_0.CLK_IN 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.2618f
C631 3bit_freq_divider_0.dff_nclk_0.nCLK a_52924_21129# 0.03449f
C632 a_64383_23628# a_64419_23326# 0.04304f
C633 a_53445_23726# a_53065_23691# 0.41048f
C634 a_54400_43159# a_54494_43159# 0.42277f
C635 a_53022_43738# a_57178_43159# 0.04095f
C636 a_51685_23725# PFD_0.VDD 0.30547f
C637 3bit_freq_divider_1.A2 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ 0.04365f
C638 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 0.02712f
C639 3bit_freq_divider_0.dff_nclk_0.D 3bit_freq_divider_0.dff_nclk_0.nRST 0.76289f
C640 a_61394_23732# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.37259f
C641 a_51600_24907# 3bit_freq_divider_0.dff_nclk_0.nRST 0.01267f
C642 PFD_0.VDD a_63426_22886# 0.20834f
C643 a_53899_22244# a_53738_22270# 0.66077f
C644 3bit_freq_divider_0.EN charge_pump_0.bias_p 0.33628f
C645 3bit_freq_divider_1.sg13g2_or3_1_0.B a_63426_22886# 0.10697f
C646 a_62654_23727# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.29516f
C647 3bit_freq_divider_0.dff_nclk_0.nCLK a_53445_23726# 0.24213f
C648 3bit_freq_divider_1.A2 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 0.15836f
C649 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_0.Cout 0.42266f
C650 m1_16847_2260# m2_16847_2260# 0.2063p
C651 a_52950_20401# PFD_0.VDD 0.2331f
C652 PFD_0.Ref_CLK PFD_0.DOWN 0.06328f
C653 PFD_0.VDD 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ 0.18067f
C654 a_53152_43159# a_52944_43077# 0.31786f
C655 a_55836_43159# a_57084_43159# 0.09682f
C656 a_64383_23889# a_64383_23706# 0.41048f
C657 3bit_freq_divider_1.freq_div_cell_0.Cin a_61878_22886# 0.01011f
C658 a_55345_24897# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.30546f
C659 3bit_freq_divider_0.EN 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.12799f
C660 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.05067f
C661 PFD_0.VDD 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 1.4225f
C662 a_60385_24947# a_60385_24717# 0.10864f
C663 3bit_freq_divider_0.dff_nclk_0.nCLK a_54504_20259# 0.37259f
C664 a_51648_21103# 3bit_freq_divider_0.sg13g2_or3_1_0.B 0.26158f
C665 sg13g2_inv_1_0.A charge_pump_0.bias_p 0.0229f
C666 PFD_0.VDD charge_pump_0.bias_p 2.67087f
C667 a_64731_24890# PFD_0.VDD 0.04155f
C668 a_54472_21129# a_54434_21392# 0.36535f
C669 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.sg13g2_or3_1_0.B 0.58488f
C670 a_53738_24026# PFD_0.VDD 0.22151f
C671 a_60967_24990# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI 0.21784f
C672 3bit_freq_divider_0.dff_nclk_0.nCLK a_53899_20488# 0.17248f
C673 a_61887_20534# a_62900_20179# 0.04306f
C674 a_59614_43129# 3bit_freq_divider_0.CLK_IN 0.09257f
C675 PFD_0.VDD a_61394_20220# 0.36995f
C676 11Stage_vco_new_0.vctl a_53147_40413# 0.04423f
C677 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 0.42892f
C678 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_60967_23234# 0.30546f
C679 a_53968_23946# PFD_0.VDD 0.32286f
C680 a_51685_23725# 3bit_freq_divider_0.A0 0.02143f
C681 3bit_freq_divider_0.EN 3bit_freq_divider_0.freq_div_cell_1.Cout 0.01552f
C682 3bit_freq_divider_0.dff_nclk_0.nCLK a_54504_22015# 0.37259f
C683 a_53774_21934# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.33731f
C684 11Stage_vco_new_0.vctl a_54627_42591# 0.07714f
C685 3bit_freq_divider_1.sg13g2_or3_1_0.C PFD_0.VDD 0.19202f
C686 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VDD 0.27798f
C687 3bit_freq_divider_1.sg13g2_nand2_1_0.Y PFD_0.VDD 3.38844f
C688 3bit_freq_divider_1.A1 m3_17285_2698# 0.2919f
C689 3bit_freq_divider_1.sg13g2_or3_1_0.C 3bit_freq_divider_1.sg13g2_or3_1_0.B 1.00414f
C690 a_53147_40413# PFD_0.VDD 0.81606f
C691 a_61887_24046# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.18489f
C692 a_63426_21130# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 0.01011f
C693 a_54627_42591# PFD_0.VDD 0.01625f
C694 charge_pump_0.bias_n charge_pump_0.bias_p 1.09436f
C695 a_63255_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 0.12248f
C696 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 0.22983f
C697 a_57111_40283# a_57173_40413# 0.1148f
C698 a_53445_23726# a_53738_24026# 0.04306f
C699 PFD_0.VDD a_60967_23234# 0.45855f
C700 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_63426_24642# 0.02246f
C701 a_51684_22284# a_51684_22692# 0.47248f
C702 3bit_freq_divider_1.dff_nclk_0.nCLK a_62900_20179# 0.2629f
C703 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.40308f
C704 a_53085_40283# a_54489_40413# 0.01208f
C705 a_63255_23244# 3bit_freq_divider_1.A2 0.01433f
C706 a_54427_40283# a_53147_40413# 0.45292f
C707 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01369f
C708 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_1.Cout 0.4595f
C709 a_54472_21129# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 0.02559f
C710 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_0.freq_div_cell_0.Cout 0.084f
C711 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.29872f
C712 3bit_freq_divider_1.dff_nclk_0.nRST a_64398_24796# 0.10221f
C713 a_61691_20534# a_61394_20220# 0.17766f
C714 a_62900_23691# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 0.10118f
C715 a_54434_24904# 3bit_freq_divider_0.freq_div_cell_0.Cin 0.01154f
C716 a_61394_21976# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 0.3562f
C717 a_62270_20543# a_62119_20605# 0.70262f
C718 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61394_20220# 0.08213f
C719 a_45451_28860# PFD_0.VDD 0.05543f
C720 3bit_freq_divider_1.CLK_OUT m6_17427_2840# 1.19758f
C721 3bit_freq_divider_1.dff_nclk_0.nRST a_64424_22200# 0.34882f
C722 a_63463_23728# PFD_0.VDD 0.2349f
C723 a_63255_23244# a_63223_22886# 0.0104f
C724 3bit_freq_divider_0.A2 3bit_freq_divider_0.EN 0.11756f
C725 a_61707_21488# PFD_0.VDD 0.2676f
C726 a_63255_23244# PFD_0.VDD 0.25835f
C727 3bit_freq_divider_0.freq_div_cell_0.Cin PFD_0.VDD 1.21627f
C728 3bit_freq_divider_0.dff_nclk_0.nCLK a_52886_21392# 0.10313f
C729 PFD_0.VDD 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 0.97883f
C730 a_63255_23244# 3bit_freq_divider_1.sg13g2_or3_1_0.B 0.23215f
C731 m3_17285_2698# m4_17285_2698# 0.20496p
C732 a_51648_24438# 3bit_freq_divider_0.dff_nclk_0.nRST 0.04054f
C733 a_53774_21934# a_53899_22244# 0.04304f
C734 a_59614_43129# PFD_0.VDD 0.44048f
C735 3bit_freq_divider_0.EN 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.02119f
C736 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.10521f
C737 a_61691_24046# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 0.01446f
C738 a_54472_24641# a_54434_24904# 0.36535f
C739 a_54504_20259# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.08213f
C740 a_53774_20178# a_53445_20214# 0.04324f
C741 a_52944_43077# PFD_0.VDD 0.88486f
C742 3bit_freq_divider_0.sg13g2_or3_1_0.C PFD_0.VDD 0.20391f
C743 a_51622_24863# a_51759_25014# 0.14868f
C744 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_1.dff_nclk_0.nCLK 0.0844f
C745 a_54472_24641# PFD_0.VDD 0.214f
C746 3bit_freq_divider_1.freq_div_cell_0.Cin a_61707_23244# 0.12082f
C747 3bit_freq_divider_1.A0 3bit_freq_divider_1.A2 0.0326f
C748 3bit_freq_divider_1.sg13g2_or3_1_0.C a_64419_23326# 0.01089f
C749 a_64383_23889# PFD_0.VDD 0.41974f
C750 a_55948_56737# 3bit_freq_divider_0.EN 0.0294f
C751 a_60584_24580# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI 0.12404f
C752 3bit_freq_divider_0.A2 PFD_0.VDD 0.25402f
C753 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.10701f
C754 a_62270_24055# a_62119_24117# 0.70262f
C755 a_51622_24863# PFD_0.VDD 0.09559f
C756 PFD_0.VDD a_53899_22244# 0.26052f
C757 PFD_0.VCO_CLK a_45658_27900# 0.17296f
C758 a_64383_23889# 3bit_freq_divider_1.dff_nclk_0.D 0.09445f
C759 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_61878_22886# 0.02559f
C760 a_51600_24907# a_51759_25014# 0.01952f
C761 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.9437f
C762 a_52924_22885# PFD_0.VDD 0.20953f
C763 3bit_freq_divider_1.A0 PFD_0.VDD 0.55412f
C764 a_64383_23628# 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.33833f
C765 a_60967_24990# 3bit_freq_divider_1.freq_div_cell_0.Cin 0.13167f
C766 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 3bit_freq_divider_1.A2 0.04535f
C767 a_56742_53480# charge_pump_0.bias_p 0.04781f
C768 a_51684_22284# a_51631_22774# 0.17766f
C769 a_51685_23725# a_51648_24041# 0.41048f
C770 a_51685_23725# a_51684_22692# 0.04306f
C771 a_53022_43738# a_55769_40283# 0.19112f
C772 a_62270_24055# PFD_0.VDD 0.26494f
C773 3bit_freq_divider_0.A2 a_52924_21129# 0.02265f
C774 a_51648_21103# a_51708_21413# 0.014f
C775 3bit_freq_divider_0.dff_nclk_0.D PFD_0.VDD 0.84532f
C776 a_64384_21091# 3bit_freq_divider_1.sg13g2_or3_1_0.A 0.31317f
C777 a_63223_21130# a_63255_21488# 0.0104f
C778 a_55831_40413# a_57112_40850# 0.22994f
C779 a_53022_43738# a_55831_40413# 0.05603f
C780 a_51600_24907# PFD_0.VDD 0.04155f
C781 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_52886_23148# 0.12248f
C782 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 1.0402f
C783 m5_17331_2744# m6_17427_2840# 84.0579f
C784 3bit_freq_divider_0.A1 a_51684_22284# 0.0269f
C785 a_55948_56737# PFD_0.VDD 0.31573f
C786 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_0.A1 0.01869f
C787 a_51693_23426# a_51684_22284# 0.45825f
C788 a_55345_21385# 3bit_freq_divider_0.freq_div_cell_1.Cout 0.13166f
C789 a_53058_43159# a_53152_43159# 0.42606f
C790 a_53022_43738# a_54494_43159# 0.0496f
C791 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ PFD_0.VDD 0.18204f
C792 a_54504_22015# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.08213f
C793 PFD_0.VDD a_61878_22886# 0.21321f
C794 PFD_0.Ref_CLK PFD_0.UP 0.15472f
C795 a_55742_43159# PFD_0.VDD 1.36686f
C796 3bit_freq_divider_0.sg13g2_or3_1_0.C 3bit_freq_divider_0.A0 0.41386f
C797 a_57178_43159# a_57311_42591# 0.22378f
C798 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_61878_24642# 0.02559f
C799 a_64459_24995# a_64398_24796# 0.0229f
C800 a_61691_24046# a_62900_23691# 0.04324f
C801 a_52944_43077# a_53285_42591# 0.03206f
C802 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_63255_25000# 0.14987f
C803 3bit_freq_divider_0.sg13g2_or3_1_0.C 3bit_freq_divider_0.sg13g2_or3_1_0.B 1.00414f
C804 a_62654_23727# a_63463_23728# 0.09575f
C805 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_54434_23148# 0.46099f
C806 a_53085_40283# PFD_0.VDD 1.35257f
C807 a_54357_49278# charge_pump_0.bias_p 0.01013f
C808 PFD_0.VDD a_51708_21299# 0.01263f
C809 a_55345_24897# 3bit_freq_divider_0.freq_div_cell_0.Cin 0.13167f
C810 a_55862_56737# charge_pump_0.bias_p 0.3307f
C811 a_54504_20259# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.3562f
C812 3bit_freq_divider_0.A2 3bit_freq_divider_0.sg13g2_or3_1_0.B 0.33008f
C813 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.02712f
C814 a_64383_23889# a_64419_23326# 0.03957f
C815 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_52950_20401# 0.12389f
C816 a_53065_20179# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ 0.0571f
C817 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.A1 0.26228f
C818 11Stage_vco_new_0.vctl a_60528_49446# 0.01545f
C819 3bit_freq_divider_0.dff_nclk_0.D 3bit_freq_divider_0.A0 0.1238f
C820 a_52924_24641# PFD_0.VDD 0.21522f
C821 3bit_freq_divider_1.freq_div_cell_1.Cout 3bit_freq_divider_0.EN 0.01552f
C822 3bit_freq_divider_0.sg13g2_or3_1_0.B a_52924_22885# 0.10697f
C823 a_61887_20534# a_62654_20215# 0.40027f
C824 a_46817_27899# PFD_0.VDD 1.02029f
C825 a_58520_43159# a_59614_43129# 0.02041f
C826 PFD_0.Ref_CLK m6_17427_2840# 1.23795f
C827 3bit_freq_divider_0.freq_div_cell_0.Cin 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 0.14552f
C828 a_51685_23725# a_51631_22774# 0.04324f
C829 a_64383_23434# 3bit_freq_divider_1.dff_nclk_0.nRST 0.126f
C830 PFD_0.VDD a_52886_24904# 0.28115f
C831 3bit_freq_divider_0.freq_div_cell_1.Cout a_54434_21392# 0.01154f
C832 a_64383_23434# a_64424_22200# 0.47248f
C833 a_54472_21129# 3bit_freq_divider_0.freq_div_cell_0.Cout 0.01011f
C834 PFD_0.VDD 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.3071f
C835 a_59799_40285# PFD_0.VDD 1.38295f
C836 a_53065_23691# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ 0.05822f
C837 a_54434_23148# a_54898_22885# 0.0104f
C838 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D a_54472_22885# 0.12185f
C839 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 0.21745f
C840 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ 0.02712f
C841 3bit_freq_divider_1.A1 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 0.15164f
C842 a_61691_24046# a_62119_24117# 0.05314f
C843 a_54472_24641# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 0.01011f
C844 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_61707_23244# 0.46099f
C845 a_53968_20434# PFD_0.VDD 0.2982f
C846 a_53774_23690# a_54504_23771# 0.17766f
C847 3bit_freq_divider_1.freq_div_cell_1.Cout PFD_0.VDD 0.4595f
C848 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ 0.02505f
C849 3bit_freq_divider_0.dff_nclk_0.nCLK a_53445_20214# 0.26292f
C850 a_62654_23727# a_62270_24055# 0.03957f
C851 3bit_freq_divider_1.dff_nclk_0.nCLK a_62654_20215# 0.31114f
C852 a_61675_21130# a_61707_21488# 0.0104f
C853 a_61887_22290# a_62900_21935# 0.04306f
C854 3bit_freq_divider_0.EN a_59097_54704# 0.03561f
C855 a_53738_22270# a_53968_22190# 0.13068f
C856 3bit_freq_divider_1.A1 3bit_freq_divider_1.A2 2.64011f
C857 a_52886_21392# a_53350_21129# 0.0104f
C858 a_51693_23075# 3bit_freq_divider_0.dff_nclk_0.nRST 0.16442f
C859 a_53065_20179# a_53738_20514# 0.40027f
C860 a_62270_22299# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.17328f
C861 a_46817_27899# a_47954_28913# 0.22374f
C862 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_55345_23141# 0.30546f
C863 a_64384_24445# a_64383_23889# 0.09575f
C864 11Stage_vco_new_0.vctl a_58454_40850# 0.04998f
C865 a_62654_23727# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 0.05822f
C866 a_61691_24046# PFD_0.VDD 0.69635f
C867 a_52924_24641# 3bit_freq_divider_0.A0 0.02265f
C868 a_52886_21392# 3bit_freq_divider_0.A2 0.39847f
C869 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ a_53445_21970# 0.10118f
C870 11Stage_vco_new_0.vctl a_53086_40850# 0.04284f
C871 a_51648_24438# PFD_0.VDD 0.24104f
C872 3bit_freq_divider_1.CLK_OUT m5_17331_2744# 0.40842f
C873 PFD_0.UP a_53147_40413# 0.01107f
C874 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_52950_22157# 0.12389f
C875 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_1.sg13g2_or3_1_0.C 0.05745f
C876 charge_pump_0.vout charge_pump_0.bias_p 0.02402f
C877 3bit_freq_divider_1.A1 PFD_0.VDD 0.44908f
C878 a_56039_25022# PFD_0.VDD 0.01215f
C879 a_53058_43159# PFD_0.VDD 1.37421f
C880 PFD_0.VDD a_61707_23244# 0.2676f
C881 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_1.Cout 0.2223f
C882 3bit_freq_divider_1.A1 3bit_freq_divider_1.sg13g2_or3_1_0.B 0.13266f
C883 3bit_freq_divider_0.sg13g2_or3_1_0.C a_51684_22692# 0.03556f
C884 PFD_0.Ref_CLK a_46749_30782# 0.97391f
C885 a_52886_24904# 3bit_freq_divider_0.A0 0.40762f
C886 3bit_freq_divider_1.sg13g2_or3_1_0.C 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.28129f
C887 3bit_freq_divider_1.dff_nclk_0.nRST a_64383_23706# 0.25925f
C888 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.dff_nclk_0.nRST 0.16209f
C889 a_54434_21392# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.24715f
C890 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.60301f
C891 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI 0.14552f
C892 a_57084_43159# PFD_0.VDD 1.35049f
C893 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_53065_21935# 0.01984f
C894 a_55769_40283# a_55831_40413# 0.12228f
C895 a_60967_24990# PFD_0.VDD 0.4548f
C896 PFD_0.VDD a_60967_21478# 0.45855f
C897 a_54504_20259# a_53968_20434# 0.45825f
C898 a_61691_22290# a_62900_21935# 0.04324f
C899 3bit_freq_divider_1.dff_nclk_0.nCLK a_61887_20534# 0.18209f
C900 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_0.Cout 0.32366f
C901 a_61887_24046# a_62270_24055# 0.66077f
C902 m7_16847_2260# 3bit_freq_divider_0.A0 1.44946f
C903 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_63463_23728# 0.12519f
C904 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D a_61878_21130# 0.12185f
C905 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.40308f
C906 a_51648_24041# 3bit_freq_divider_0.dff_nclk_0.D 0.09445f
C907 3bit_freq_divider_0.dff_nclk_0.D a_51684_22692# 0.0175f
C908 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ a_63463_20216# 0.21609f
C909 a_55836_43159# a_55969_42591# 0.22378f
C910 a_47777_29803# PFD_0.VDD 1.07957f
C911 a_53968_20434# a_53899_20488# 0.70262f
C912 a_53065_21935# a_53445_21970# 0.41048f
C913 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ a_52950_22157# 0.21609f
C914 a_61394_23732# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.08213f
C915 a_51648_24438# 3bit_freq_divider_0.A0 0.01187f
C916 a_64383_23300# 3bit_freq_divider_1.dff_nclk_0.nRST 0.31482f
C917 a_59097_54704# charge_pump_0.bias_n 0.01331f
C918 a_58536_54976# charge_pump_0.bias_p 0.38944f
C919 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_0.A2 0.17317f
C920 a_64383_23300# a_64424_22200# 0.45825f
C921 a_55862_56737# a_55948_56737# 0.0609f
C922 a_52944_43077# PFD_0.UP 0.01107f
C923 a_54489_40413# a_55770_40850# 0.2342f
C924 a_53022_43738# a_53147_40413# 0.10922f
C925 a_53445_21970# a_53738_22270# 0.04306f
C926 a_54842_49733# PFD_0.VDD 0.03367f
C927 3bit_freq_divider_0.dff_nclk_0.nCLK a_53774_20178# 0.35517f
C928 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.22983f
C929 a_60479_25023# PFD_0.VDD 0.01215f
C930 a_62654_21971# a_62900_21935# 0.41048f
C931 a_63463_21972# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.05956f
C932 a_59799_40285# a_58520_43159# 0.12666f
C933 a_53065_21935# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ 0.0571f
C934 PFD_0.VDD a_63463_20216# 0.2331f
C935 a_53350_24641# a_52886_24904# 0.0104f
C936 a_61691_24046# a_61394_23732# 0.17766f
C937 a_64362_24865# a_64731_24890# 0.01952f
C938 PFD_0.VDD 3bit_freq_divider_0.sg13g2_or3_1_0.A 0.12791f
C939 11Stage_vco_new_0.vctl a_57173_40413# 0.02576f
C940 a_61691_24046# a_62654_23727# 0.02302f
C941 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.40308f
C942 a_53774_21934# a_53968_22190# 0.05314f
C943 a_53065_23691# a_53899_24000# 0.03957f
C944 a_53738_24026# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01324f
C945 a_54747_49259# PFD_0.DOWN 0.01456f
C946 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 3bit_freq_divider_1.dff_nclk_0.nCLK 0.21745f
C947 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_1.A0 0.20944f
C948 a_63426_24642# a_63255_25000# 0.36535f
C949 3bit_freq_divider_0.sg13g2_or3_1_0.C 3bit_freq_divider_0.A1 0.20623f
C950 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ PFD_0.VDD 0.18065f
C951 a_57173_40413# PFD_0.VDD 1.11589f
C952 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_62654_20215# 0.01984f
C953 3bit_freq_divider_0.A0 m4_17285_2698# 0.39515f
C954 3bit_freq_divider_0.dff_nclk_0.nCLK a_53899_24000# 0.17312f
C955 a_53065_21935# a_52950_22157# 0.09575f
C956 a_61878_21130# 3bit_freq_divider_1.freq_div_cell_0.Cout 0.01011f
C957 3bit_freq_divider_0.A2 3bit_freq_divider_0.A1 0.01072f
C958 3bit_freq_divider_0.sg13g2_or3_1_0.A a_52924_21129# 0.10614f
C959 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.60301f
C960 a_58520_43159# a_58454_40850# 0.02056f
C961 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 0.02712f
C962 a_52886_23148# a_53350_22885# 0.0104f
C963 a_56887_49467# a_56695_49467# 0.01287f
C964 a_61887_24046# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01324f
C965 a_64384_21091# PFD_0.VDD 0.34084f
C966 3bit_freq_divider_0.A1 a_52924_22885# 0.02265f
C967 a_64384_21091# 3bit_freq_divider_1.sg13g2_or3_1_0.B 0.26158f
C968 3bit_freq_divider_0.dff_nclk_0.D a_51631_22774# 0.03728f
C969 a_60584_24580# PFD_0.VDD 0.10495f
C970 PFD_0.VDD a_53968_22190# 0.31854f
C971 a_64398_24796# PFD_0.VDD 0.09559f
C972 a_61691_22290# a_61887_22290# 0.45047f
C973 PFD_0.Ref_CLK m5_17331_2744# 0.42278f
C974 3bit_freq_divider_0.sg13g2_nand2_1_0.Y a_55345_23141# 0.08797f
C975 a_53022_43738# a_52944_43077# 0.97477f
C976 a_56887_49467# charge_pump_0.vout 0.63953f
C977 PFD_0.VDD a_62119_20605# 0.2982f
C978 3bit_freq_divider_1.dff_nclk_0.nRST PFD_0.VDD 0.60883f
C979 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_0.Cin 0.084f
C980 PFD_0.VDD a_62270_20543# 0.24492f
C981 3bit_freq_divider_0.dff_nclk_0.D 3bit_freq_divider_0.A1 0.11556f
C982 PFD_0.VDD a_64424_22200# 0.36995f
C983 a_56828_53480# sg13g2_inv_1_0.A 0.06208f
C984 3bit_freq_divider_0.dff_nclk_0.D a_51693_23426# 0.04146f
C985 3bit_freq_divider_1.A0 m6_17427_2840# 1.19758f
C986 a_53065_23691# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.02071f
C987 3bit_freq_divider_1.dff_nclk_0.nRST 3bit_freq_divider_1.dff_nclk_0.D 0.7629f
C988 m1_17285_2698# 3bit_freq_divider_0.A0 0.01061f
C989 a_57111_40283# PFD_0.VDD 1.36202f
C990 3bit_freq_divider_1.dff_nclk_0.D a_64424_22200# 0.43097f
C991 11Stage_vco_new_0.vctl a_55836_43159# 0.02165f
C992 a_61878_21130# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 0.02559f
C993 a_53065_21935# a_53738_22270# 0.40027f
C994 a_62900_21935# 3bit_freq_divider_1.A2 0.0145f
C995 a_52886_23148# PFD_0.VDD 0.25998f
C996 a_61691_24046# a_61887_24046# 0.45047f
C997 a_51693_23075# PFD_0.VDD 0.2446f
C998 a_53738_20514# PFD_0.VDD 0.19386f
C999 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.08441f
C1000 3bit_freq_divider_0.freq_div_cell_0.Cin 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01369f
C1001 a_64383_23434# a_64383_23706# 0.04306f
C1002 3bit_freq_divider_0.sg13g2_or3_1_0.B 3bit_freq_divider_0.sg13g2_or3_1_0.A 0.72102f
C1003 a_63255_21488# 3bit_freq_divider_1.sg13g2_or3_1_0.A 0.23182f
C1004 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_0.Cout 0.32366f
C1005 3bit_freq_divider_0.freq_div_cell_1.Cout 3bit_freq_divider_0.freq_div_cell_0.Cout 0.09134f
C1006 a_55836_43159# PFD_0.VDD 1.18255f
C1007 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_53774_20178# 0.33731f
C1008 a_51648_24041# a_51648_24438# 0.09575f
C1009 3bit_freq_divider_0.freq_div_cell_0.Cout 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01369f
C1010 a_61887_22290# a_62654_21971# 0.40027f
C1011 3bit_freq_divider_0.EN a_58734_56203# 0.07729f
C1012 a_59799_40285# a_58515_40413# 0.45428f
C1013 a_45658_27900# a_46817_27899# 0.43194f
C1014 3bit_freq_divider_1.dff_nclk_0.nCLK a_63426_22886# 0.03415f
C1015 11Stage_vco_new_0.vctl a_55770_40850# 0.05041f
C1016 a_62900_21935# PFD_0.VDD 0.30801f
C1017 a_53774_21934# a_53445_21970# 0.04324f
C1018 a_53738_24026# a_53899_24000# 0.66077f
C1019 3bit_freq_divider_0.freq_div_cell_0.Cin 3bit_freq_divider_0.freq_div_cell_0.Cout 0.10559f
C1020 11Stage_vco_new_0.vctl a_58653_42591# 0.08336f
C1021 a_61691_20534# a_62119_20605# 0.05314f
C1022 a_56038_24617# PFD_0.VDD 0.0448f
C1023 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.22983f
C1024 a_61691_20534# a_62270_20543# 0.04304f
C1025 a_61394_20220# a_61887_20534# 0.47248f
C1026 PFD_0.VDD 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI 0.7718f
C1027 a_56828_53480# charge_pump_0.bias_n 0.01798f
C1028 a_61675_22886# a_61707_23244# 0.0104f
C1029 a_53022_43738# a_55742_43159# 0.19603f
C1030 PFD_0.VDD a_55770_40850# 0.01475f
C1031 3bit_freq_divider_1.sg13g2_or3_1_0.C a_63426_24642# 0.10662f
C1032 PFD_0.VDD a_54434_23148# 0.2676f
C1033 a_63463_21972# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ 0.21609f
C1034 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q PFD_0.VDD 1.42273f
C1035 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ 0.0874f
C1036 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VDD 0.28742f
C1037 a_53968_23946# a_53899_24000# 0.70262f
C1038 3bit_freq_divider_0.dff_nclk_0.nCLK a_53065_23691# 0.29533f
C1039 a_53774_23690# PFD_0.VDD 0.70098f
C1040 3bit_freq_divider_0.dff_nclk_0.nCLK a_51648_21103# 0.33244f
C1041 3bit_freq_divider_1.A2 3bit_freq_divider_1.sg13g2_or3_1_0.A 0.10441f
C1042 a_64383_23300# a_64383_23434# 0.13068f
C1043 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.freq_div_cell_0.Cout 0.01369f
C1044 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 1.04018f
C1045 a_60528_49446# charge_pump_0.vout 0.01545f
C1046 PFD_0.VDD a_58734_56203# 0.35557f
C1047 a_61707_25000# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI 0.12082f
C1048 a_58515_40413# a_58454_40850# 0.03282f
C1049 a_53022_43738# a_53085_40283# 0.2302f
C1050 3bit_freq_divider_1.dff_nclk_0.nRST a_64419_23326# 0.16457f
C1051 PFD_0.VDD a_53445_21970# 0.30838f
C1052 a_54504_20259# a_53738_20514# 0.47248f
C1053 a_54504_22015# a_53968_22190# 0.45825f
C1054 PFD_0.VDD 3bit_freq_divider_1.sg13g2_or3_1_0.A 0.12797f
C1055 3bit_freq_divider_1.sg13g2_or3_1_0.A 3bit_freq_divider_1.sg13g2_or3_1_0.B 0.72102f
C1056 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 0.22983f
C1057 3bit_freq_divider_1.dff_nclk_0.nCLK a_61394_20220# 0.37259f
C1058 a_61691_22290# a_62654_21971# 0.02302f
C1059 a_61707_21488# a_61878_21130# 0.36535f
C1060 a_52886_21392# 3bit_freq_divider_0.sg13g2_or3_1_0.A 0.23182f
C1061 a_52886_23148# 3bit_freq_divider_0.sg13g2_or3_1_0.B 0.23215f
C1062 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 0.21603f
C1063 3bit_freq_divider_1.A1 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 0.18013f
C1064 a_53738_20514# a_53899_20488# 0.66077f
C1065 a_64459_24995# PFD_0.VDD 0.08543f
C1066 a_53445_23726# a_53774_23690# 0.04324f
C1067 a_54494_43159# a_54627_42591# 0.22417f
C1068 a_45579_29803# PFD_0.VDD 0.45874f
C1069 3bit_freq_divider_1.sg13g2_or3_1_0.C 3bit_freq_divider_1.dff_nclk_0.nCLK 0.13894f
C1070 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_1.dff_nclk_0.nCLK 0.23907f
C1071 a_54504_23771# PFD_0.VDD 0.38531f
C1072 PFD_0.VDD 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ 0.18275f
C1073 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D a_61394_20220# 0.3562f
C1074 a_53147_40413# a_54428_40850# 0.2377f
C1075 a_53022_43738# a_59799_40285# 0.19389f
C1076 3bit_freq_divider_0.dff_nclk_0.nCLK a_52950_20401# 0.05883f
C1077 a_53774_20178# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.01446f
C1078 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.05067f
C1079 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_60967_24990# 0.30546f
C1080 a_61394_21976# a_61887_22290# 0.47248f
C1081 a_63426_21130# 3bit_freq_divider_1.sg13g2_or3_1_0.A 0.10614f
C1082 PFD_0.VDD a_55345_23141# 0.45855f
C1083 a_53065_21935# a_53774_21934# 0.02335f
C1084 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.CLK_IN 0.2618f
C1085 m6_17427_2840# m7_16847_2260# 25.5177f
C1086 a_53738_24026# a_53065_23691# 0.40027f
C1087 PFD_0.VDD a_56137_24678# 0.11858f
C1088 a_61887_22290# PFD_0.VDD 0.21577f
C1089 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 0.42266f
C1090 m7_16847_2260# PFD_0.VSS 93.0612f
C1091 m6_17427_2840# PFD_0.VSS 0.10708p
C1092 m6_16847_2260# PFD_0.VSS 0.11472p
C1093 m5_17331_2744# PFD_0.VSS 79.2024f
C1094 m5_16847_2260# PFD_0.VSS 84.4749f
C1095 m4_17285_2698# PFD_0.VSS 84.41901f
C1096 m4_16847_2260# PFD_0.VSS 89.24989f
C1097 m3_17285_2698# PFD_0.VSS 91.8291f
C1098 m3_16847_2260# PFD_0.VSS 96.21301f
C1099 m2_17285_2698# PFD_0.VSS 0.10557p
C1100 m2_16847_2260# PFD_0.VSS 0.10679p
C1101 m1_17285_2698# PFD_0.VSS 0.22685p
C1102 m1_16847_2260# PFD_0.VSS 0.22893p
C1103 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ PFD_0.VSS 0.08893f $ **FLOATING
C1104 a_62900_20179# PFD_0.VSS 0.34783f $ **FLOATING
C1105 a_63463_20216# PFD_0.VSS 0.43565f $ **FLOATING
C1106 a_62654_20215# PFD_0.VSS 0.80634f $ **FLOATING
C1107 a_62119_20605# PFD_0.VSS 0.26895f $ **FLOATING
C1108 a_62270_20543# PFD_0.VSS 0.16883f $ **FLOATING
C1109 a_61887_20534# PFD_0.VSS 1.05953f $ **FLOATING
C1110 a_61394_20220# PFD_0.VSS 0.13262f $ **FLOATING
C1111 a_61691_20534# PFD_0.VSS 0.79964f $ **FLOATING
C1112 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VSS 0.51487f $ **FLOATING
C1113 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VSS 0.51489f $ **FLOATING
C1114 a_54504_20259# PFD_0.VSS 0.13262f $ **FLOATING
C1115 a_53899_20488# PFD_0.VSS 0.16883f $ **FLOATING
C1116 a_53968_20434# PFD_0.VSS 0.26896f $ **FLOATING
C1117 a_53738_20514# PFD_0.VSS 1.05953f $ **FLOATING
C1118 a_53445_20214# PFD_0.VSS 0.34783f $ **FLOATING
C1119 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ PFD_0.VSS 0.08893f $ **FLOATING
C1120 a_53774_20178# PFD_0.VSS 0.80054f $ **FLOATING
C1121 a_53065_20179# PFD_0.VSS 0.80634f $ **FLOATING
C1122 a_52950_20401# PFD_0.VSS 0.43566f $ **FLOATING
C1123 a_64384_21091# PFD_0.VSS 0.59054f $ **FLOATING
C1124 3bit_freq_divider_1.sg13g2_or3_1_0.A PFD_0.VSS 0.77543f $ **FLOATING
C1125 a_63255_21488# PFD_0.VSS 0.38381f $ **FLOATING
C1126 3bit_freq_divider_1.A2 PFD_0.VSS 0.12039p $ **FLOATING
C1127 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D PFD_0.VSS 0.49782f $ **FLOATING
C1128 a_61707_21488# PFD_0.VSS 0.36496f $ **FLOATING
C1129 3bit_freq_divider_1.freq_div_cell_1.Cout PFD_0.VSS 0.14556f $ **FLOATING
C1130 a_60967_21478# PFD_0.VSS 0.27989f $ **FLOATING
C1131 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q PFD_0.VSS 2.25165f $ **FLOATING
C1132 3bit_freq_divider_0.freq_div_cell_1.Cout PFD_0.VSS 0.14556f $ **FLOATING
C1133 a_55345_21385# PFD_0.VSS 0.27989f $ **FLOATING
C1134 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D PFD_0.VSS 0.49784f $ **FLOATING
C1135 a_54434_21392# PFD_0.VSS 0.36496f $ **FLOATING
C1136 3bit_freq_divider_0.sg13g2_or3_1_0.A PFD_0.VSS 0.77447f $ **FLOATING
C1137 a_51648_21103# PFD_0.VSS 0.59026f $ **FLOATING
C1138 3bit_freq_divider_0.A2 PFD_0.VSS 91.68561f $ **FLOATING
C1139 a_52886_21392# PFD_0.VSS 0.3838f $ **FLOATING
C1140 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q PFD_0.VSS 2.25169f $ **FLOATING
C1141 a_60922_21796# PFD_0.VSS 0.03012f $ **FLOATING
C1142 a_60922_21818# PFD_0.VSS 0.02768f $ **FLOATING
C1143 a_52808_21795# PFD_0.VSS 0.03012f $ **FLOATING
C1144 a_52808_21817# PFD_0.VSS 0.02768f $ **FLOATING
C1145 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VSS 0.50854f $ **FLOATING
C1146 a_64424_22200# PFD_0.VSS 0.12168f $ **FLOATING
C1147 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ PFD_0.VSS 0.07921f $ **FLOATING
C1148 a_62900_21935# PFD_0.VSS 0.33549f $ **FLOATING
C1149 a_63463_21972# PFD_0.VSS 0.42316f $ **FLOATING
C1150 a_62654_21971# PFD_0.VSS 0.7639f $ **FLOATING
C1151 a_62119_22361# PFD_0.VSS 0.25006f $ **FLOATING
C1152 a_62270_22299# PFD_0.VSS 0.1501f $ **FLOATING
C1153 a_61887_22290# PFD_0.VSS 1.02135f $ **FLOATING
C1154 a_61394_21976# PFD_0.VSS 0.12168f $ **FLOATING
C1155 a_61691_22290# PFD_0.VSS 0.77938f $ **FLOATING
C1156 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VSS 0.47143f $ **FLOATING
C1157 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VSS 0.47143f $ **FLOATING
C1158 a_54504_22015# PFD_0.VSS 0.12168f $ **FLOATING
C1159 a_53899_22244# PFD_0.VSS 0.1501f $ **FLOATING
C1160 a_53968_22190# PFD_0.VSS 0.25006f $ **FLOATING
C1161 a_53738_22270# PFD_0.VSS 1.02135f $ **FLOATING
C1162 a_53445_21970# PFD_0.VSS 0.33549f $ **FLOATING
C1163 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ PFD_0.VSS 0.07921f $ **FLOATING
C1164 a_53774_21934# PFD_0.VSS 0.78026f $ **FLOATING
C1165 a_53065_21935# PFD_0.VSS 0.7639f $ **FLOATING
C1166 a_52950_22157# PFD_0.VSS 0.4233f $ **FLOATING
C1167 3bit_freq_divider_1.sg13g2_or3_1_0.B PFD_0.VSS 1.39257f $ **FLOATING
C1168 a_64383_23300# PFD_0.VSS 0.25093f $ **FLOATING
C1169 a_63255_23244# PFD_0.VSS 0.37914f $ **FLOATING
C1170 3bit_freq_divider_1.A1 PFD_0.VSS 0.10102p $ **FLOATING
C1171 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D PFD_0.VSS 0.45601f $ **FLOATING
C1172 a_61707_23244# PFD_0.VSS 0.36159f $ **FLOATING
C1173 3bit_freq_divider_1.freq_div_cell_0.Cout PFD_0.VSS 1.80113f $ **FLOATING
C1174 a_60967_23234# PFD_0.VSS 0.27786f $ **FLOATING
C1175 a_64419_23326# PFD_0.VSS 0.1501f $ **FLOATING
C1176 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q PFD_0.VSS 2.24178f $ **FLOATING
C1177 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VSS 0.50854f $ **FLOATING
C1178 a_51684_22284# PFD_0.VSS 0.12168f $ **FLOATING
C1179 3bit_freq_divider_0.freq_div_cell_0.Cout PFD_0.VSS 1.80115f $ **FLOATING
C1180 a_55345_23141# PFD_0.VSS 0.27786f $ **FLOATING
C1181 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D PFD_0.VSS 0.45601f $ **FLOATING
C1182 a_54434_23148# PFD_0.VSS 0.36159f $ **FLOATING
C1183 3bit_freq_divider_0.sg13g2_or3_1_0.B PFD_0.VSS 1.39146f $ **FLOATING
C1184 3bit_freq_divider_0.A1 PFD_0.VSS 94.7177f $ **FLOATING
C1185 a_52886_23148# PFD_0.VSS 0.37912f $ **FLOATING
C1186 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q PFD_0.VSS 2.2418f $ **FLOATING
C1187 a_64383_23628# PFD_0.VSS 0.82074f $ **FLOATING
C1188 a_64383_23434# PFD_0.VSS 1.02665f $ **FLOATING
C1189 a_60922_23552# PFD_0.VSS 0.03012f $ **FLOATING
C1190 a_60922_23574# PFD_0.VSS 0.02768f $ **FLOATING
C1191 a_52808_23551# PFD_0.VSS 0.03012f $ **FLOATING
C1192 a_52808_23573# PFD_0.VSS 0.02768f $ **FLOATING
C1193 a_51693_23426# PFD_0.VSS 0.25093f $ **FLOATING
C1194 a_51693_23075# PFD_0.VSS 0.1501f $ **FLOATING
C1195 a_64383_23706# PFD_0.VSS 0.33666f $ **FLOATING
C1196 3bit_freq_divider_1.dff_nclk_0.D PFD_0.VSS 0.57206f $ **FLOATING
C1197 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ PFD_0.VSS 0.08281f $ **FLOATING
C1198 a_62900_23691# PFD_0.VSS 0.33612f $ **FLOATING
C1199 a_63463_23728# PFD_0.VSS 0.42235f $ **FLOATING
C1200 a_62654_23727# PFD_0.VSS 0.76426f $ **FLOATING
C1201 a_62119_24117# PFD_0.VSS 0.25006f $ **FLOATING
C1202 a_62270_24055# PFD_0.VSS 0.1501f $ **FLOATING
C1203 a_61887_24046# PFD_0.VSS 1.02191f $ **FLOATING
C1204 a_61394_23732# PFD_0.VSS 0.12168f $ **FLOATING
C1205 a_61691_24046# PFD_0.VSS 0.78738f $ **FLOATING
C1206 3bit_freq_divider_1.dff_nclk_0.nCLK PFD_0.VSS 7.48134f $ **FLOATING
C1207 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VSS 0.47246f $ **FLOATING
C1208 a_51631_22774# PFD_0.VSS 0.82147f $ **FLOATING
C1209 a_51684_22692# PFD_0.VSS 1.02713f $ **FLOATING
C1210 3bit_freq_divider_1.sg13g2_nand2_1_0.Y PFD_0.VSS 2.56526f $ **FLOATING
C1211 3bit_freq_divider_0.sg13g2_nand2_1_0.Y PFD_0.VSS 2.56527f $ **FLOATING
C1212 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK PFD_0.VSS 0.47246f $ **FLOATING
C1213 a_54504_23771# PFD_0.VSS 0.12168f $ **FLOATING
C1214 a_53899_24000# PFD_0.VSS 0.1501f $ **FLOATING
C1215 a_53968_23946# PFD_0.VSS 0.25006f $ **FLOATING
C1216 a_53738_24026# PFD_0.VSS 1.02191f $ **FLOATING
C1217 a_53445_23726# PFD_0.VSS 0.33612f $ **FLOATING
C1218 3bit_freq_divider_0.dff_nclk_0.nCLK PFD_0.VSS 7.50548f $ **FLOATING
C1219 a_51685_23725# PFD_0.VSS 0.33666f $ **FLOATING
C1220 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ PFD_0.VSS 0.08281f $ **FLOATING
C1221 a_53774_23690# PFD_0.VSS 0.78853f $ **FLOATING
C1222 a_53065_23691# PFD_0.VSS 0.76426f $ **FLOATING
C1223 a_52950_23913# PFD_0.VSS 0.42231f $ **FLOATING
C1224 a_64383_23889# PFD_0.VSS 0.79267f $ **FLOATING
C1225 a_64384_24445# PFD_0.VSS 0.41218f $ **FLOATING
C1226 3bit_freq_divider_1.CLK_OUT PFD_0.VSS 92.2343f $ **FLOATING
C1227 3bit_freq_divider_0.dff_nclk_0.D PFD_0.VSS 0.57206f $ **FLOATING
C1228 a_51648_24041# PFD_0.VSS 0.7928f $ **FLOATING
C1229 3bit_freq_divider_1.dff_nclk_0.nRST PFD_0.VSS 1.21235f $ **FLOATING
C1230 a_64398_24796# PFD_0.VSS 0.17085f $ **FLOATING
C1231 a_64338_24910# PFD_0.VSS 0.01158f $ **FLOATING
C1232 a_64362_24865# PFD_0.VSS 0.18902f $ **FLOATING
C1233 a_64459_24995# PFD_0.VSS 0.21807f $ **FLOATING
C1234 a_51648_24438# PFD_0.VSS 0.41218f $ **FLOATING
C1235 3bit_freq_divider_1.sg13g2_or3_1_0.C PFD_0.VSS 2.00849f $ **FLOATING
C1236 a_63255_25000# PFD_0.VSS 0.38174f $ **FLOATING
C1237 3bit_freq_divider_1.A0 PFD_0.VSS 92.142f $ **FLOATING
C1238 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D PFD_0.VSS 0.4595f $ **FLOATING
C1239 a_61707_25000# PFD_0.VSS 0.36409f $ **FLOATING
C1240 3bit_freq_divider_1.freq_div_cell_0.Cin PFD_0.VSS 1.81006f $ **FLOATING
C1241 a_60967_24990# PFD_0.VSS 0.27856f $ **FLOATING
C1242 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q PFD_0.VSS 2.27033f $ **FLOATING
C1243 a_60584_24580# PFD_0.VSS 0.16608f $ **FLOATING
C1244 a_60385_24947# PFD_0.VSS 0.21087f $ **FLOATING
C1245 a_56137_24678# PFD_0.VSS 0.21087f $ **FLOATING
C1246 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI PFD_0.VSS 1.60229f $ **FLOATING
C1247 a_60385_24717# PFD_0.VSS 0.17977f $ **FLOATING
C1248 a_60479_25023# PFD_0.VSS 0.01118f $ **FLOATING
C1249 a_55941_24882# PFD_0.VSS 0.16608f $ **FLOATING
C1250 3bit_freq_divider_0.dff_nclk_0.nRST PFD_0.VSS 1.20799f $ **FLOATING
C1251 a_51622_24863# PFD_0.VSS 0.17085f $ **FLOATING
C1252 3bit_freq_divider_0.freq_div_cell_0.Cin PFD_0.VSS 1.81006f $ **FLOATING
C1253 a_55345_24897# PFD_0.VSS 0.27856f $ **FLOATING
C1254 a_56039_25022# PFD_0.VSS 0.01118f $ **FLOATING
C1255 a_56013_24979# PFD_0.VSS 0.17977f $ **FLOATING
C1256 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D PFD_0.VSS 0.4595f $ **FLOATING
C1257 a_54434_24904# PFD_0.VSS 0.36409f $ **FLOATING
C1258 3bit_freq_divider_0.sg13g2_or3_1_0.C PFD_0.VSS 2.00844f $ **FLOATING
C1259 a_52065_24890# PFD_0.VSS 0.01158f $ **FLOATING
C1260 a_51721_24988# PFD_0.VSS 0.21807f $ **FLOATING
C1261 a_51759_25014# PFD_0.VSS 0.18902f $ **FLOATING
C1262 3bit_freq_divider_0.A0 PFD_0.VSS 90.2415f $ **FLOATING
C1263 a_52886_24904# PFD_0.VSS 0.38144f $ **FLOATING
C1264 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI PFD_0.VSS 1.60229f $ **FLOATING
C1265 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q PFD_0.VSS 2.27033f $ **FLOATING
C1266 a_47954_28913# PFD_0.VSS 0.97627f $ **FLOATING
C1267 a_46817_27899# PFD_0.VSS 1.26528f $ **FLOATING
C1268 a_45658_27900# PFD_0.VSS 1.24513f $ **FLOATING
C1269 PFD_0.VCO_CLK PFD_0.VSS 5.09845f $ **FLOATING
C1270 a_48909_28913# PFD_0.VSS 1.03223f $ **FLOATING
C1271 a_45451_28860# PFD_0.VSS 1.00878f $ **FLOATING
C1272 a_47777_29803# PFD_0.VSS 1.2524f $ **FLOATING
C1273 a_46749_30782# PFD_0.VSS 1.31435f $ **FLOATING
C1274 a_45579_29803# PFD_0.VSS 0.97532f $ **FLOATING
C1275 PFD_0.Ref_CLK PFD_0.VSS 93.6639f $ **FLOATING
C1276 a_59799_40285# PFD_0.VSS 0.05405f $ **FLOATING
C1277 a_58453_40283# PFD_0.VSS 0.0472f $ **FLOATING
C1278 a_57111_40283# PFD_0.VSS 0.04799f $ **FLOATING
C1279 a_55769_40283# PFD_0.VSS 0.04714f $ **FLOATING
C1280 a_54427_40283# PFD_0.VSS 0.0482f $ **FLOATING
C1281 a_53085_40283# PFD_0.VSS 0.0663f $ **FLOATING
C1282 a_58515_40413# PFD_0.VSS 5.02759f $ **FLOATING
C1283 a_57173_40413# PFD_0.VSS 5.13846f $ **FLOATING
C1284 a_55831_40413# PFD_0.VSS 5.22541f $ **FLOATING
C1285 a_54489_40413# PFD_0.VSS 5.4642f $ **FLOATING
C1286 a_53147_40413# PFD_0.VSS 5.81185f $ **FLOATING
C1287 a_59800_40852# PFD_0.VSS 0.75356f $ **FLOATING
C1288 a_58454_40850# PFD_0.VSS 0.80499f $ **FLOATING
C1289 a_57112_40850# PFD_0.VSS 0.81838f $ **FLOATING
C1290 a_55770_40850# PFD_0.VSS 0.83004f $ **FLOATING
C1291 a_54428_40850# PFD_0.VSS 0.82862f $ **FLOATING
C1292 a_53086_40850# PFD_0.VSS 0.83267f $ **FLOATING
C1293 a_59600_42432# PFD_0.VSS 0.27494f $ **FLOATING
C1294 a_58653_42591# PFD_0.VSS 0.65274f $ **FLOATING
C1295 a_57311_42591# PFD_0.VSS 0.67166f $ **FLOATING
C1296 a_55969_42591# PFD_0.VSS 0.67176f $ **FLOATING
C1297 a_54627_42591# PFD_0.VSS 0.67671f $ **FLOATING
C1298 a_53285_42591# PFD_0.VSS 0.68456f $ **FLOATING
C1299 3bit_freq_divider_0.CLK_IN PFD_0.VSS 22.1194f $ **FLOATING
C1300 a_59614_43129# PFD_0.VSS 0.26077f $ **FLOATING
C1301 a_58520_43159# PFD_0.VSS 6.8154f $ **FLOATING
C1302 a_57178_43159# PFD_0.VSS 5.12501f $ **FLOATING
C1303 a_55836_43159# PFD_0.VSS 4.87283f $ **FLOATING
C1304 a_54494_43159# PFD_0.VSS 4.85892f $ **FLOATING
C1305 a_53152_43159# PFD_0.VSS 5.07652f $ **FLOATING
C1306 a_52944_43077# PFD_0.VSS 5.94106f $ **FLOATING
C1307 a_58426_43159# PFD_0.VSS 0.05881f $ **FLOATING
C1308 a_57084_43159# PFD_0.VSS 0.03948f $ **FLOATING
C1309 a_55742_43159# PFD_0.VSS 0.04155f $ **FLOATING
C1310 a_54400_43159# PFD_0.VSS 0.04203f $ **FLOATING
C1311 a_53058_43159# PFD_0.VSS 0.05441f $ **FLOATING
C1312 a_53022_43738# PFD_0.VSS 5.38922f $ **FLOATING
C1313 a_54747_49259# PFD_0.VSS 0.16684f $ **FLOATING
C1314 PFD_0.DOWN PFD_0.VSS 13.9137f $ **FLOATING
C1315 a_60528_49446# PFD_0.VSS 0.16044f
C1316 a_56695_49467# PFD_0.VSS 0.14015f
C1317 11Stage_vco_new_0.vctl PFD_0.VSS 17.2488f $ **FLOATING
C1318 a_56887_49467# PFD_0.VSS 8.04158f $ **FLOATING
C1319 a_54357_49278# PFD_0.VSS 0.26592f $ **FLOATING
C1320 PFD_0.UP PFD_0.VSS 12.6584f $ **FLOATING
C1321 charge_pump_0.vout PFD_0.VSS 28.7608f $ **FLOATING
C1322 a_56828_53480# PFD_0.VSS 2.32258f
C1323 a_56742_53480# PFD_0.VSS 1.67237f $ **FLOATING
C1324 a_59097_54704# PFD_0.VSS 0.1681f $ **FLOATING
C1325 a_58536_54976# PFD_0.VSS 0.61525f $ **FLOATING
C1326 a_58734_56203# PFD_0.VSS 0.05948f $ **FLOATING
C1327 charge_pump_0.bias_p PFD_0.VSS 5.47872f $ **FLOATING
C1328 charge_pump_0.bias_n PFD_0.VSS 6.55127f $ **FLOATING
C1329 3bit_freq_divider_0.EN PFD_0.VSS 51.6717f $ **FLOATING
C1330 sg13g2_inv_1_0.A PFD_0.VSS 0.10244p $ **FLOATING
C1331 a_55948_56737# PFD_0.VSS 1.95792f
C1332 a_55862_56737# PFD_0.VSS 0.99714f $ **FLOATING
C1333 PFD_0.VDD PFD_0.VSS 0.19478p $ **FLOATING
.ends
