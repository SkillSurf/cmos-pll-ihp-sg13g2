* Extracted by KLayout with SG13G2 LVS runset on : 10/06/2025 18:11

.SUBCKT t2_or4
M$1 4 3 5 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u PD=0.74u
M$2 5 3 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u PD=1.34u
M$3 6 4 7 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u PD=0.74u
M$4 7 9 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u PD=1.34u
M$5 9 8 10 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$6 10 8 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$7 11 6 12 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$8 12 6 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$9 13 11 14 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$10 14 15 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$11 15 16 17 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$12 17 16 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$13 19 18 20 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$14 20 18 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$15 16 19 21 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$16 21 23 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$17 23 22 24 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$18 24 22 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$19 1 3 4 1 sg13_lv_pmos L=0.13u W=0.6u AS=0.159p AD=0.159p PS=1.96u PD=1.96u
M$21 1 4 6 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$22 6 9 1 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$23 1 8 9 1 sg13_lv_pmos L=0.13u W=0.6u AS=0.159p AD=0.159p PS=1.96u PD=1.96u
M$25 1 6 11 1 sg13_lv_pmos L=0.13u W=0.6u AS=0.159p AD=0.159p PS=1.96u PD=1.96u
M$27 1 11 13 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$28 13 15 1 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$29 1 16 15 1 sg13_lv_pmos L=0.13u W=0.6u AS=0.159p AD=0.159p PS=1.96u PD=1.96u
M$31 1 18 19 1 sg13_lv_pmos L=0.13u W=0.6u AS=0.159p AD=0.159p PS=1.96u PD=1.96u
M$33 1 19 16 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$34 16 23 1 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$35 1 22 23 1 sg13_lv_pmos L=0.13u W=0.6u AS=0.159p AD=0.159p PS=1.96u PD=1.96u
.ENDS t2_or4
