** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_dff_2_tb.sch
**.subckt t2_dff_2_tb
Vs VDD GND 1.2
* noconn Q
* noconn QN
Vdin D GND dc 0 ac 0 pulse(0, 1.2, 0, 50p, 50p, 2.5n, 5n)
Vclk CLK GND dc 0 ac 0 pulse(0, 1.2, 0, 50p, 50p, 1.25n, 2.5n)
Vrst RST GND dc 0 ac 0 pulse(0, 1.2, 0, 50p, 50p, 8n, 15n)
x1 D CLK Q VDD QN RST GND t2_dff_2
**** begin user architecture code


.param temp=27
.control
save all
tran 10p 15n
write tran_t2_dff_2.raw
.endc



.lib cornerMOSlv.lib mos_ff

**** end user architecture code
**.ends

* expanding   symbol:  t2_dff_2.sym # of pins=7
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_dff_2.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_dff_2.sch
.subckt t2_dff_2 D nCLK Q VDD nQ nRST VSS
*.iopin VSS
*.ipin D
*.ipin nRST
*.opin Q
*.iopin VDD
*.opin nQ
*.ipin nCLK
XM1 net1 D VDD VDD sg13_lv_pmos w=0.3u l=0.15u ng=1 m=1
XM2 net2 CLK net1 VDD sg13_lv_pmos w=0.3u l=0.15u ng=1 m=1
XM3 net2 D VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM4 net3 CLK VDD VDD sg13_lv_pmos w=0.3u l=0.15u ng=1 m=1
XM6 net4 CLK VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM5 net3 net2 net4 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM7 nQ net3 VDD VDD sg13_lv_pmos w=0.3u l=0.15u ng=1 m=1
XM8 net5 net3 VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM9 nQ CLK net5 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM10 nQ nRST VDD VDD sg13_lv_pmos w=0.3u l=0.15u ng=1 m=1
XM11 Q nQ VDD VDD sg13_lv_pmos w=0.3u l=0.15u ng=1 m=1
XM12 Q nQ VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
x1 VDD nCLK CLK VSS t2_inverter
.ends


* expanding   symbol:  t2_inverter.sym # of pins=4
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_inverter.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_inverter.sch
.subckt t2_inverter VP A Y VN
*.iopin VP
*.iopin VN
*.ipin A
*.opin Y
XM2 Y A VP VP sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
XM1 Y A VN VN sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
