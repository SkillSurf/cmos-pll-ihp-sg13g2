** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_bias.sch
.subckt t2_bias VPWR VPB VGND VNB en bias_n bias_p enb
*.PININFO VPWR:B VPB:B VGND:B VNB:B en:I enb:I bias_n:O bias_p:O
M9 net1 en VPWR VPB sg13_lv_pmos w=0.5u l=0.15u ng=1 m=1
M10 bias_p bias_p VPWR VPB sg13_lv_pmos w=0.2u l=1.0u ng=1 m=5
M1 dio_mid dio_mid VPWR VPB sg13_lv_pmos w=0.5u l=0.15u ng=1 m=1
M2 net1 net1 dio_mid VPB sg13_lv_pmos w=0.5u l=0.15u ng=1 m=1
M3 bias_p en VPWR VPB sg13_lv_pmos w=0.5u l=0.15u ng=1 m=1
M4 bias_n bias_p res_bot VPB sg13_lv_pmos w=0.2u l=1.0u ng=1 m=5
M11 kick_sw en VGND VNB sg13_lv_nmos w=0.5u l=0.15u ng=1 m=1
M12 bias_p net1 kick_sw VNB sg13_lv_nmos w=0.5u l=0.15u ng=1 m=1
M5 net1 bias_n VGND VNB sg13_lv_nmos w=0.2u l=1.0u ng=1 m=5
M6 bias_p bias_n VGND VNB sg13_lv_nmos w=0.2u l=1.0u ng=1 m=5
M7 bias_n enb VGND VNB sg13_lv_nmos w=0.5u l=0.15u ng=1 m=1
M8 bias_n bias_n VGND VNB sg13_lv_nmos w=0.2u l=1.0u ng=1 m=5
R1 res_bot VPWR rhigh w=0.5e-6 l=0.5e-6 m=1 b=0
.ends
