** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_or4.sch
.subckt t2_or4 VDD VSS inA inB inC inD out
*.PININFO VSS:B inD:I out:O VDD:B inA:I inB:I inC:I
x1 VDD VSS inA inB net2 t2_or2
x2 VDD VSS inC inD net1 t2_or2
x3 VDD VSS net2 net1 out t2_or2
.ends

* expanding   symbol:  t2_or2.sym # of pins=5
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_or2.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_or2.sch
.subckt t2_or2 VDD VSS inA inB out
*.PININFO VSS:B inA:I inB:I out:O VDD:B
x2 VDD inA inA net2 VSS t2_nand2
x3 VDD inB inB net1 VSS t2_nand2
x4 VDD net2 net1 out VSS t2_nand2
.ends


* expanding   symbol:  t2_nand2.sym # of pins=5
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand2.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand2.sch
.subckt t2_nand2 VDD inA inB out VSS
*.PININFO VSS:B inA:I inB:I out:O VDD:B
M1 out inA VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M2 out inB VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M3 out inB net1 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M4 net1 inA VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends

