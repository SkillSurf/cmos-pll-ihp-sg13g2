.subckt 11Stage_vco_new_update2 VDD VSS
.ends
.end
