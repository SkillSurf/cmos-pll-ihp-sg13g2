** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/charge_pump.sch
.subckt charge_pump VP bias_p up vout down bias_n VN
*.PININFO bias_p:I up:I down:I bias_n:I VN:B VP:B vout:O
M1 net1 bias_n VN VN sg13_lv_nmos w=1.2u l=0.13u ng=1 m=1
M2 vout down net1 VN sg13_lv_nmos w=1.2u l=0.13u ng=1 m=1
M3 vout net3 net2 VP sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
M4 net2 bias_p VP VP sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
x1 VP up net3 VN inverter
.ends

* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /foss/designs/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/inverter.sym
** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/inverter.sch
.subckt inverter VP IN OUT VN
*.PININFO VN:B VP:B IN:I OUT:O
M1 OUT IN VN VN sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M2 OUT IN VP VP sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
.ends

