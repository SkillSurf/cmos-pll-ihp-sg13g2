* Extracted by KLayout with SG13G2 LVS runset on : 10/07/2025 15:19

.SUBCKT 11Stage_vco_new
M$1 \$85 \$47 \$54 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$2 \$54 \$47 \$85 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p
+ PS=0.74u PD=1.34u
M$3 \$86 \$48 \$47 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$4 \$47 \$48 \$86 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p
+ PS=0.74u PD=1.34u
M$5 \$87 \$49 \$48 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$6 \$48 \$49 \$87 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p
+ PS=0.74u PD=1.34u
M$7 \$88 \$50 \$49 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$8 \$49 \$50 \$88 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p
+ PS=0.74u PD=1.34u
M$9 \$89 \$51 \$50 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$10 \$50 \$51 \$89 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p
+ PS=0.74u PD=1.34u
M$11 \$90 \$52 \$51 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$12 \$51 \$52 \$90 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p
+ PS=0.74u PD=1.34u
M$13 \$106 \$104 \$85 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p
+ PS=1.28u PD=0.74u
M$14 \$85 \$104 \$106 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p
+ PS=0.74u PD=1.28u
M$15 \$107 \$104 \$86 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p
+ PS=1.28u PD=0.74u
M$16 \$86 \$104 \$107 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p
+ PS=0.74u PD=1.28u
M$17 \$108 \$104 \$87 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p
+ PS=1.28u PD=0.74u
M$18 \$87 \$104 \$108 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p
+ PS=0.74u PD=1.28u
M$19 \$109 \$104 \$88 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p
+ PS=1.28u PD=0.74u
M$20 \$88 \$104 \$109 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p
+ PS=0.74u PD=1.28u
M$21 \$110 \$104 \$89 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p
+ PS=1.28u PD=0.74u
M$22 \$89 \$104 \$110 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p
+ PS=0.74u PD=1.28u
M$23 \$1 \$104 \$11 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p
+ PS=1.28u PD=0.74u
M$24 \$11 \$104 \$1 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p
+ PS=0.74u PD=1.28u
M$25 \$124 \$104 \$125 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p
+ PS=1.28u PD=0.74u
M$26 \$125 \$104 \$124 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p
+ PS=0.74u PD=1.28u
M$27 \$126 \$104 \$127 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p
+ PS=1.28u PD=0.74u
M$28 \$127 \$104 \$126 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p
+ PS=0.74u PD=1.28u
M$29 \$128 \$104 \$129 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p
+ PS=1.28u PD=0.74u
M$30 \$129 \$104 \$128 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p
+ PS=0.74u PD=1.28u
M$31 \$130 \$104 \$131 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p
+ PS=1.28u PD=0.74u
M$32 \$131 \$104 \$130 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p
+ PS=0.74u PD=1.28u
M$33 \$132 \$104 \$133 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p
+ PS=1.28u PD=0.74u
M$34 \$133 \$104 \$132 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p
+ PS=0.74u PD=1.28u
M$35 \$111 \$104 \$90 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p
+ PS=1.28u PD=0.74u
M$36 \$90 \$104 \$111 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p
+ PS=0.74u PD=1.28u
M$37 \$125 \$54 \$146 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$38 \$146 \$54 \$125 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p
+ PS=0.74u PD=1.34u
M$39 \$127 \$146 \$147 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$40 \$147 \$146 \$127 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p
+ PS=0.74u PD=1.34u
M$41 \$129 \$147 \$148 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$42 \$148 \$147 \$129 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p
+ PS=0.74u PD=1.34u
M$43 \$131 \$148 \$149 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$44 \$149 \$148 \$131 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p
+ PS=0.74u PD=1.34u
M$45 \$133 \$149 \$52 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$46 \$52 \$149 \$133 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p
+ PS=0.74u PD=1.34u
M$47 \$1 \$52 \$37 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$48 \$37 \$52 \$1 \$1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p
+ PS=0.74u PD=1.34u
M$49 \$6 \$11 \$4 \$41 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p
+ PS=0.745u PD=1.34u
M$50 \$4 \$11 \$6 \$41 sg13_lv_pmos L=0.13u W=0.2u AS=0.104p AD=0.059p PS=1.34u
+ PD=0.74u
M$51 \$6 \$11 \$4 \$41 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u
+ PD=0.74u
M$52 \$6 \$11 \$4 \$41 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p
+ PS=0.745u PD=0.74u
M$53 \$7 \$11 \$4 \$42 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p
+ PS=0.745u PD=1.34u
M$54 \$4 \$11 \$7 \$42 sg13_lv_pmos L=0.13u W=0.2u AS=0.104p AD=0.059p PS=1.34u
+ PD=0.74u
M$55 \$7 \$11 \$4 \$42 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u
+ PD=0.74u
M$56 \$7 \$11 \$4 \$42 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p
+ PS=0.745u PD=0.74u
M$57 \$8 \$11 \$4 \$44 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p
+ PS=0.745u PD=1.34u
M$58 \$4 \$11 \$8 \$44 sg13_lv_pmos L=0.13u W=0.2u AS=0.104p AD=0.059p PS=1.34u
+ PD=0.74u
M$59 \$8 \$11 \$4 \$44 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u
+ PD=0.74u
M$60 \$8 \$11 \$4 \$44 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p
+ PS=0.745u PD=0.74u
M$61 \$9 \$11 \$4 \$46 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p
+ PS=0.745u PD=1.34u
M$62 \$4 \$11 \$9 \$46 sg13_lv_pmos L=0.13u W=0.2u AS=0.104p AD=0.059p PS=1.34u
+ PD=0.74u
M$63 \$9 \$11 \$4 \$46 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u
+ PD=0.74u
M$64 \$9 \$11 \$4 \$46 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p
+ PS=0.745u PD=0.74u
M$65 \$10 \$11 \$4 \$45 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p
+ PS=0.745u PD=1.34u
M$66 \$4 \$11 \$10 \$45 sg13_lv_pmos L=0.13u W=0.2u AS=0.104p AD=0.059p
+ PS=1.34u PD=0.74u
M$67 \$10 \$11 \$4 \$45 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p
+ PS=0.74u PD=0.74u
M$68 \$10 \$11 \$4 \$45 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p
+ PS=0.745u PD=0.74u
M$69 \$54 \$47 \$6 \$80 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.1075p
+ PS=0.745u PD=1.34u
M$70 \$6 \$47 \$54 \$80 sg13_lv_pmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$71 \$54 \$47 \$6 \$80 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.0625p
+ PS=0.74u PD=0.74u
M$72 \$54 \$47 \$6 \$80 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.0625p
+ PS=0.745u PD=0.74u
M$73 \$47 \$48 \$7 \$82 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.1075p
+ PS=0.745u PD=1.34u
M$74 \$7 \$48 \$47 \$82 sg13_lv_pmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$75 \$47 \$48 \$7 \$82 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.0625p
+ PS=0.74u PD=0.74u
M$76 \$47 \$48 \$7 \$82 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.0625p
+ PS=0.745u PD=0.74u
M$77 \$48 \$49 \$8 \$84 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.1075p
+ PS=0.745u PD=1.34u
M$78 \$8 \$49 \$48 \$84 sg13_lv_pmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$79 \$48 \$49 \$8 \$84 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.0625p
+ PS=0.74u PD=0.74u
M$80 \$48 \$49 \$8 \$84 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.0625p
+ PS=0.745u PD=0.74u
M$81 \$49 \$50 \$9 \$83 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.1075p
+ PS=0.745u PD=1.34u
M$82 \$9 \$50 \$49 \$83 sg13_lv_pmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$83 \$49 \$50 \$9 \$83 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.0625p
+ PS=0.74u PD=0.74u
M$84 \$49 \$50 \$9 \$83 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.0625p
+ PS=0.745u PD=0.74u
M$85 \$50 \$51 \$10 \$81 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.1075p
+ PS=0.745u PD=1.34u
M$86 \$10 \$51 \$50 \$81 sg13_lv_pmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$87 \$50 \$51 \$10 \$81 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.0625p
+ PS=0.74u PD=0.74u
M$88 \$50 \$51 \$10 \$81 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.0625p
+ PS=0.745u PD=0.74u
M$89 \$12 \$11 \$4 \$43 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p
+ PS=0.745u PD=1.34u
M$90 \$4 \$11 \$12 \$43 sg13_lv_pmos L=0.13u W=0.2u AS=0.104p AD=0.059p
+ PS=1.34u PD=0.74u
M$91 \$12 \$11 \$4 \$43 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p
+ PS=0.74u PD=0.74u
M$92 \$12 \$11 \$4 \$43 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p
+ PS=0.745u PD=0.74u
M$93 \$4 \$11 \$11 \$5 sg13_lv_pmos L=0.13u W=0.2u AS=0.104p AD=0.059p PS=1.34u
+ PD=0.74u
M$94 \$11 \$11 \$4 \$5 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u
+ PD=0.74u
M$95 \$4 \$11 \$11 \$5 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.05975p
+ PS=0.74u PD=0.745u
M$96 \$11 \$11 \$4 \$5 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p
+ PS=0.745u PD=1.34u
M$97 \$146 \$54 \$161 \$174 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.0625p
+ PS=0.745u PD=0.74u
M$98 \$161 \$54 \$146 \$174 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.0625p
+ PS=0.74u PD=0.74u
M$99 \$146 \$54 \$161 \$174 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p
+ PS=0.74u PD=1.34u
M$100 \$146 \$54 \$161 \$174 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p
+ AD=0.1075p PS=0.745u PD=1.34u
M$101 \$147 \$146 \$162 \$179 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p
+ AD=0.0625p PS=0.745u PD=0.74u
M$102 \$162 \$146 \$147 \$179 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p
+ AD=0.0625p PS=0.74u PD=0.74u
M$103 \$147 \$146 \$162 \$179 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p
+ AD=0.1075p PS=0.74u PD=1.34u
M$104 \$147 \$146 \$162 \$179 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p
+ AD=0.1075p PS=0.745u PD=1.34u
M$105 \$148 \$147 \$163 \$184 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p
+ AD=0.0625p PS=0.745u PD=0.74u
M$106 \$163 \$147 \$148 \$184 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p
+ AD=0.0625p PS=0.74u PD=0.74u
M$107 \$148 \$147 \$163 \$184 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p
+ AD=0.1075p PS=0.74u PD=1.34u
M$108 \$148 \$147 \$163 \$184 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p
+ AD=0.1075p PS=0.745u PD=1.34u
M$109 \$149 \$148 \$164 \$191 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p
+ AD=0.0625p PS=0.745u PD=0.74u
M$110 \$164 \$148 \$149 \$191 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p
+ AD=0.0625p PS=0.74u PD=0.74u
M$111 \$149 \$148 \$164 \$191 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p
+ AD=0.1075p PS=0.74u PD=1.34u
M$112 \$149 \$148 \$164 \$191 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p
+ AD=0.1075p PS=0.745u PD=1.34u
M$113 \$52 \$149 \$165 \$192 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p
+ AD=0.0625p PS=0.745u PD=0.74u
M$114 \$165 \$149 \$52 \$192 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.0625p
+ PS=0.74u PD=0.74u
M$115 \$52 \$149 \$165 \$192 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p
+ PS=0.74u PD=1.34u
M$116 \$52 \$149 \$165 \$192 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p
+ AD=0.1075p PS=0.745u PD=1.34u
M$117 \$51 \$52 \$12 \$79 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.1075p
+ PS=0.745u PD=1.34u
M$118 \$12 \$52 \$51 \$79 sg13_lv_pmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p
+ PS=1.34u PD=0.74u
M$119 \$51 \$52 \$12 \$79 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.0625p
+ PS=0.74u PD=0.74u
M$120 \$51 \$52 \$12 \$79 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.0625p
+ PS=0.745u PD=0.74u
M$121 \$4 \$52 \$37 \$160 sg13_lv_pmos L=0.13u W=0.2u AS=0.104p AD=0.059p
+ PS=1.34u PD=0.74u
M$122 \$37 \$52 \$4 \$160 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p
+ PS=0.74u PD=0.74u
M$123 \$4 \$52 \$166 \$160 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p
+ PS=0.74u PD=0.74u
M$124 \$166 \$52 \$4 \$160 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.104p
+ PS=0.74u PD=1.34u
M$125 \$161 \$11 \$4 \$202 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p
+ PS=0.745u PD=0.74u
M$126 \$4 \$11 \$196 \$202 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p
+ PS=0.74u PD=0.74u
M$127 \$196 \$11 \$4 \$202 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.104p
+ PS=0.74u PD=1.34u
M$128 \$161 \$11 \$4 \$202 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p
+ PS=0.745u PD=1.34u
M$129 \$162 \$11 \$4 \$207 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p
+ PS=0.745u PD=0.74u
M$130 \$4 \$11 \$162 \$207 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p
+ PS=0.74u PD=0.74u
M$131 \$162 \$11 \$4 \$207 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.104p
+ PS=0.74u PD=1.34u
M$132 \$162 \$11 \$4 \$207 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p
+ PS=0.745u PD=1.34u
M$133 \$163 \$11 \$4 \$212 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p
+ PS=0.745u PD=0.74u
M$134 \$4 \$11 \$163 \$212 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p
+ PS=0.74u PD=0.74u
M$135 \$163 \$11 \$4 \$212 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.104p
+ PS=0.74u PD=1.34u
M$136 \$163 \$11 \$4 \$212 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p
+ PS=0.745u PD=1.34u
M$137 \$164 \$11 \$4 \$218 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p
+ PS=0.745u PD=0.74u
M$138 \$4 \$11 \$164 \$218 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p
+ PS=0.74u PD=0.74u
M$139 \$164 \$11 \$4 \$218 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.104p
+ PS=0.74u PD=1.34u
M$140 \$164 \$11 \$4 \$218 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p
+ PS=0.745u PD=1.34u
M$141 \$165 \$11 \$4 \$213 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p
+ PS=0.745u PD=0.74u
M$142 \$4 \$11 \$165 \$213 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p
+ PS=0.74u PD=0.74u
M$143 \$165 \$11 \$4 \$213 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.104p
+ PS=0.74u PD=1.34u
M$144 \$165 \$11 \$4 \$213 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p
+ PS=0.745u PD=1.34u
C$145 \$3 \$48 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$146 \$3 \$52 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$147 \$3 \$49 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$148 \$3 \$50 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$149 \$3 \$2 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$150 \$3 \$37 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$151 \$3 \$47 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$152 \$3 \$54 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$153 \$3 \$147 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$154 \$3 \$148 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$155 \$3 \$37 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$156 \$3 \$146 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$157 \$3 \$149 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
.ENDS 11Stage_vco_new
