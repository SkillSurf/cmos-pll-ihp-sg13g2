* Extracted by KLayout with SG13G2 LVS runset on : 06/07/2025 12:18

.SUBCKT TOP
X$1 12 10 8 1 10 pmos$1
X$2 12 7 8 1 7 pmos$2
X$3 5 11 5 8 1 7 7 pmos
X$4 7 6 1 9 nmos$1
X$5 9 3 1 5 nmos$2
X$6 12 11 1 rppd
X$7 7 3 1 5 nmos$2
X$8 5 3 1 5 nmos$2
X$9 5 3 1 2 nmos$1
X$10 6 3 1 4 nmos$1
X$11 12 7 8 1 4 pmos$1
X$12 10 9 8 1 9 pmos$1
X$13 12 9 8 1 4 pmos$1
.ENDS TOP

.SUBCKT rppd 1 2 3
R$1 1 2 rppd w=1u l=4u ps=0 b=0 m=1
.ENDS rppd

.SUBCKT nmos$2 1 2 3 4
M$1 1 4 2 3 sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
.ENDS nmos$2

.SUBCKT nmos$1 1 2 3 4
M$1 1 4 2 3 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
.ENDS nmos$1

.SUBCKT pmos 1 2 3 4 5 6 7
M$1 1 6 2 4 sg13_lv_pmos L=1u W=2u AS=0.68p AD=0.38p PS=4.68u PD=2.38u
M$2 2 7 3 4 sg13_lv_pmos L=1u W=2u AS=0.38p AD=0.68p PS=2.38u PD=4.68u
.ENDS pmos

.SUBCKT pmos$2 1 2 3 4 5
M$1 1 5 2 3 sg13_lv_pmos L=1u W=2u AS=0.68p AD=0.68p PS=4.68u PD=4.68u
.ENDS pmos$2

.SUBCKT pmos$1 1 2 3 4 5
M$1 1 5 2 3 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
.ENDS pmos$1
