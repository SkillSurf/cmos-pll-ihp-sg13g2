** sch_path: /foss/designs/tutorials/inverter/inverter_tb.sch
**.subckt inverter_tb
V1 VDD GND 1.2
Vin Vin GND PULSE(0 1.2 .2NS .2NS .2NS 5NS 10NS)
x1 net1 Vin net2 net3 inverter
**** begin user architecture code


.include= /foss/designs/tutorials/inverter/output_RC/inverter__inverter/magic_RC/inverter.pex.spice
.param temp=27
.tran 1p 30n uic
.save all


 .lib cornerMOSlv.lib mos_tt

**** end user architecture code
**.ends

* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /foss/designs/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/inverter.sym
** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/inverter.sch
.subckt inverter VP IN OUT VN
*.iopin VN
*.iopin VP
*.ipin IN
*.opin OUT
XM1 OUT IN VN VN sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM2 OUT IN VP VP sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
