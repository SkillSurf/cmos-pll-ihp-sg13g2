* NGSPICE file created from half_add.ext - technology: ihp-sg13g2

.subckt half_add inA sum inB VDD VSS cout
X0 VSS a_57_n6# sum VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X1 VSS inB a_n589_n14# VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.1216p ps=1.02u w=0.64u l=0.13u
X2 a_n589_n14# inA a_n683_n14# VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.2176p ps=1.96u w=0.64u l=0.13u
X3 VSS inB a_57_n6# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X4 VDD inA a_228_238# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X5 a_228_238# inB VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X6 a_57_n6# inB a_25_262# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X7 cout a_n683_n14# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1331p ps=1.12u w=0.74u l=0.13u
X8 VDD inB a_n683_n14# VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.1596p ps=1.22u w=0.84u l=0.13u
X9 sum a_57_n6# a_228_238# VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X10 a_n683_n14# inA VDD VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.2856p ps=2.36u w=0.84u l=0.13u
X11 cout a_n683_n14# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.1918p ps=1.5u w=1.12u l=0.13u
X12 a_25_262# inA VDD VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X13 a_322_n44# inA VSS VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X14 sum inB a_322_n44# VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X15 a_57_n6# inA VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
C0 a_n683_n14# inB 0.30545f
C1 sum VDD 0.08235f
C2 a_228_238# VDD 0.20834f
C3 cout VDD 0.29974f
C4 sum a_228_238# 0.11602f
C5 a_n683_n14# inA 0.13033f
C6 inB VDD 0.31435f
C7 a_57_n6# VDD 0.25468f
C8 sum inB 0.08794f
C9 a_57_n6# sum 0.24142f
C10 inB a_228_238# 0.02512f
C11 a_57_n6# a_228_238# 0.36535f
C12 inB cout 0.22229f
C13 a_57_n6# cout 0.01154f
C14 inA VDD 0.28939f
C15 a_57_n6# inB 0.45519f
C16 a_n683_n14# VDD 0.43783f
C17 a_228_238# inA 0.01011f
C18 cout inA 0.07689f
C19 a_25_262# a_57_n6# 0.0104f
C20 a_n683_n14# cout 0.13166f
C21 inB inA 0.42207f
C22 a_57_n6# inA 0.12082f
R0 VSS.n6 VSS.n5 1455.25
R1 VSS.n3 VSS.n1 17.001
R2 VSS.n1 VSS.n0 17.0005
R3 VSS.n5 VSS.n4 3.1147
R4 VSS VSS.n6 0.417695
R5 VSS.n6 VSS 0.298933
R6 VSS.n4 VSS 0.2055
R7 VSS VSS.n0 0.0605
R8 VSS.n3 VSS.n2 0.0351579
R9 VSS.n2 VSS 0.0228929
R10 VSS.n2 VSS.n0 0.01175
R11 VSS.n4 VSS.n3 0.00885683
R12 VSS.n5 VSS.n1 0.0010117
R13 inA.n4 inA.n2 9.81991
R14 inA.n2 inA.n1 9.01785
R15 inA.n4 inA.n3 7.50513
R16 inA.n1 inA.n0 7.501
R17 inA.n2 inA 0.0702658
R18 inA inA.n4 0.0654197
R19 inA.n1 inA 0.0505118
R20 inB.n4 inB.n1 15.1844
R21 inB.n6 inB.n0 15.0231
R22 inB.n3 inB.n2 15.0005
R23 inB.n6 inB.n5 10.5511
R24 inB.n5 inB.n4 9.0005
R25 inB.n5 inB 0.466263
R26 inB.n4 inB.n3 0.187664
R27 inB inB.n6 0.0625513
R28 inB.n3 inB 0.0513955
C23 sum VSS 0.30557f
C24 cout VSS 0.21277f
C25 inB VSS 1.0967f
C26 inA VSS 1.52964f
C27 VDD VSS 0.29349f
C28 a_57_n6# VSS 0.37141f $ **FLOATING
C29 a_n683_n14# VSS 0.32069f $ **FLOATING
.ends
