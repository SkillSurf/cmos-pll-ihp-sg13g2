* Extracted by KLayout with SG13G2 LVS runset on : 10/06/2025 18:06

.SUBCKT t2_xor2
M$1 4 3 5 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u PD=0.74u
M$2 5 6 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u PD=1.34u
M$3 6 3 7 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u PD=0.74u
M$4 7 10 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$5 8 4 9 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u PD=0.74u
M$6 9 11 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$7 11 6 12 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$8 12 10 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$9 1 3 4 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$10 4 6 1 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$11 1 3 6 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$12 6 10 1 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$13 1 4 8 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$14 8 11 1 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$15 1 6 11 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$16 11 10 1 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u PD=1.28u
.ENDS t2_xor2
