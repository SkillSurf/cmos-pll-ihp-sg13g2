* Extracted by KLayout with SG13G2 LVS runset on : 10/06/2025 08:09

.SUBCKT t2_nand2
M$1 \$1 \$5 \$3 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$2 \$3 \$6 \$4 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$3 \$2 \$5 \$4 \$2 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u
+ PD=0.68u
M$4 \$4 \$6 \$2 \$2 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u
+ PD=1.28u
.ENDS t2_nand2
