* Extracted by KLayout with SG13G2 LVS runset on : 23/07/2025 18:55

.SUBCKT 11Stage_vco_new VGND VPWR vctl Vout
M$1 VGND vctl \$136 VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.102 AD=0.066 PS=1.28
+ PD=0.74
M$2 \$136 vctl VGND VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.066 AD=0.102 PS=0.74
+ PD=1.28
M$3 VGND vctl \$130 VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.102 AD=0.066 PS=1.28
+ PD=0.74
M$4 \$130 vctl VGND VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.066 AD=0.102 PS=0.74
+ PD=1.28
M$5 VGND vctl \$124 VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.102 AD=0.066 PS=1.28
+ PD=0.74
M$6 \$124 vctl VGND VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.066 AD=0.102 PS=0.74
+ PD=1.28
M$7 VGND vctl \$127 VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.102 AD=0.066 PS=1.28
+ PD=0.74
M$8 \$127 vctl VGND VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.066 AD=0.102 PS=0.74
+ PD=1.28
M$9 VGND vctl \$86 VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.102 AD=0.066 PS=1.28
+ PD=0.74
M$10 \$86 vctl VGND VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.066 AD=0.102 PS=0.74
+ PD=1.28
M$11 VGND vctl \$84 VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.102 AD=0.066 PS=1.28
+ PD=0.74
M$12 \$84 vctl VGND VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.066 AD=0.102 PS=0.74
+ PD=1.28
M$13 VGND vctl \$83 VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.102 AD=0.066 PS=1.28
+ PD=0.74
M$14 \$83 vctl VGND VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.066 AD=0.102 PS=0.74
+ PD=1.28
M$15 \$84 \$64 \$44 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$16 \$44 \$64 \$84 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
M$17 \$81 \$59 \$51 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$18 \$51 \$59 \$81 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
M$19 VGND vctl \$85 VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.102 AD=0.066 PS=1.28
+ PD=0.74
M$20 \$85 vctl VGND VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.066 AD=0.102 PS=0.74
+ PD=1.28
M$21 \$86 \$45 \$40 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$22 \$40 \$45 \$86 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
M$23 \$83 \$44 \$48 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$24 \$48 \$44 \$83 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
M$25 \$85 \$40 \$64 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$26 \$64 \$40 \$85 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
M$27 VGND vctl \$125 VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.102 AD=0.066 PS=1.28
+ PD=0.74
M$28 \$125 vctl VGND VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.066 AD=0.102 PS=0.74
+ PD=1.28
M$29 \$82 \$48 \$59 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$30 \$59 \$48 \$82 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
M$31 VGND vctl \$82 VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.102 AD=0.066 PS=1.28
+ PD=0.74
M$32 \$82 vctl VGND VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.066 AD=0.102 PS=0.74
+ PD=1.28
M$33 VGND vctl \$39 VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.102 AD=0.066 PS=1.28
+ PD=0.74
M$34 \$39 vctl VGND VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.066 AD=0.102 PS=0.74
+ PD=1.28
M$35 VGND vctl \$81 VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.102 AD=0.066 PS=1.28
+ PD=0.74
M$36 \$81 vctl VGND VGND sg13_lv_nmos L=0.13 W=0.3 AS=0.066 AD=0.102 PS=0.74
+ PD=1.28
M$37 \$155 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.059
+ PS=0.745 PD=0.74
M$38 VPWR \$39 \$155 VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.059 PS=0.74
+ PD=0.74
M$39 \$155 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.104 PS=0.74
+ PD=1.34
M$40 \$155 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.104
+ PS=0.745 PD=1.34
M$41 \$152 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.059
+ PS=0.745 PD=0.74
M$42 VPWR \$39 \$152 VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.059 PS=0.74
+ PD=0.74
M$43 \$152 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.104 PS=0.74
+ PD=1.34
M$44 \$152 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.104
+ PS=0.745 PD=1.34
M$45 \$153 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.059
+ PS=0.745 PD=0.74
M$46 VPWR \$39 \$153 VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.059 PS=0.74
+ PD=0.74
M$47 \$153 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.104 PS=0.74
+ PD=1.34
M$48 \$153 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.104
+ PS=0.745 PD=1.34
M$49 \$156 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.059
+ PS=0.745 PD=0.74
M$50 VPWR \$39 \$156 VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.059 PS=0.74
+ PD=0.74
M$51 \$156 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.104 PS=0.74
+ PD=1.34
M$52 \$156 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.104
+ PS=0.745 PD=1.34
M$53 \$154 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.059
+ PS=0.745 PD=0.74
M$54 VPWR \$39 \$154 VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.059 PS=0.74
+ PD=0.74
M$55 \$154 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.104 PS=0.74
+ PD=1.34
M$56 \$154 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.104
+ PS=0.745 PD=1.34
M$57 \$40 \$45 \$8 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.17 PS=0.945
+ PD=1.68
M$58 \$8 \$45 \$40 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$59 \$40 \$45 \$8 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.11 PS=0.94
+ PD=0.94
M$60 \$40 \$45 \$8 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.11 PS=0.945
+ PD=0.94
M$61 \$64 \$40 \$7 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.17 PS=0.945
+ PD=1.68
M$62 \$7 \$40 \$64 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$63 \$64 \$40 \$7 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.11 PS=0.94
+ PD=0.94
M$64 \$64 \$40 \$7 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.11 PS=0.945
+ PD=0.94
M$65 \$4 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.104 PS=0.745
+ PD=1.34
M$66 VPWR \$39 \$4 VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.104 AD=0.059 PS=1.34
+ PD=0.74
M$67 \$4 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.059 PS=0.74
+ PD=0.74
M$68 \$4 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.059 PS=0.745
+ PD=0.74
M$69 \$8 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.104 PS=0.745
+ PD=1.34
M$70 VPWR \$39 \$8 VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.104 AD=0.059 PS=1.34
+ PD=0.74
M$71 \$8 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.059 PS=0.74
+ PD=0.74
M$72 \$8 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.059 PS=0.745
+ PD=0.74
M$73 \$5 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.104 PS=0.745
+ PD=1.34
M$74 VPWR \$39 \$5 VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.104 AD=0.059 PS=1.34
+ PD=0.74
M$75 \$5 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.059 PS=0.74
+ PD=0.74
M$76 \$5 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.059 PS=0.745
+ PD=0.74
M$77 \$44 \$64 \$6 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.17 PS=0.945
+ PD=1.68
M$78 \$6 \$64 \$44 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$79 \$44 \$64 \$6 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.11 PS=0.94
+ PD=0.94
M$80 \$44 \$64 \$6 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.11 PS=0.945
+ PD=0.94
M$81 \$7 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.104 PS=0.745
+ PD=1.34
M$82 VPWR \$39 \$7 VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.104 AD=0.059 PS=1.34
+ PD=0.74
M$83 \$7 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.059 PS=0.74
+ PD=0.74
M$84 \$7 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.059 PS=0.745
+ PD=0.74
M$85 \$6 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.104 PS=0.745
+ PD=1.34
M$86 VPWR \$39 \$6 VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.104 AD=0.059 PS=1.34
+ PD=0.74
M$87 \$6 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.059 PS=0.74
+ PD=0.74
M$88 \$6 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.059 PS=0.745
+ PD=0.74
M$89 \$59 \$48 \$4 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.17 PS=0.945
+ PD=1.68
M$90 \$4 \$48 \$59 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$91 \$59 \$48 \$4 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.11 PS=0.94
+ PD=0.94
M$92 \$59 \$48 \$4 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.11 PS=0.945
+ PD=0.94
M$93 \$51 \$59 \$3 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.17 PS=0.945
+ PD=1.68
M$94 \$3 \$59 \$51 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$95 \$51 \$59 \$3 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.11 PS=0.94
+ PD=0.94
M$96 \$51 \$59 \$3 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.11 PS=0.945
+ PD=0.94
M$97 \$48 \$44 \$5 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.17 PS=0.945
+ PD=1.68
M$98 \$5 \$44 \$48 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$99 \$48 \$44 \$5 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.11 PS=0.94
+ PD=0.94
M$100 \$48 \$44 \$5 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.11 PS=0.945
+ PD=0.94
M$101 \$3 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.104 PS=0.745
+ PD=1.34
M$102 VPWR \$39 \$3 VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.104 AD=0.059 PS=1.34
+ PD=0.74
M$103 \$3 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.059 PS=0.74
+ PD=0.74
M$104 \$3 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.059 PS=0.745
+ PD=0.74
M$105 VPWR \$39 \$39 VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.104 AD=0.059 PS=1.34
+ PD=0.74
M$106 \$39 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.059 PS=0.74
+ PD=0.74
M$107 VPWR \$39 \$39 VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.059 AD=0.05975 PS=0.74
+ PD=0.745
M$108 \$39 \$39 VPWR VPWR sg13_lv_pmos L=0.13 W=0.2 AS=0.05975 AD=0.104
+ PS=0.745 PD=1.34
M$109 VGND \$45 Vout VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$110 Vout \$45 VGND VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
M$111 VPWR \$45 Vout VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$112 Vout \$45 VPWR VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.11 PS=0.94
+ PD=0.94
M$113 VPWR \$45 Vout VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.11 PS=0.94
+ PD=0.94
M$114 Vout \$45 VPWR VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
C$115 \$48 VGND cap_cmim w=6.99 l=6.99 A=48.8601 P=27.96 m=1
C$116 Vout VGND cap_cmim w=6.99 l=6.99 A=48.8601 P=27.96 m=1
C$117 \$142 VGND cap_cmim w=6.99 l=6.99 A=48.8601 P=27.96 m=1
C$118 \$59 VGND cap_cmim w=6.99 l=6.99 A=48.8601 P=27.96 m=1
C$119 \$143 VGND cap_cmim w=6.99 l=6.99 A=48.8601 P=27.96 m=1
C$120 \$64 VGND cap_cmim w=6.99 l=6.99 A=48.8601 P=27.96 m=1
C$121 \$144 VGND cap_cmim w=6.99 l=6.99 A=48.8601 P=27.96 m=1
C$122 \$145 VGND cap_cmim w=6.99 l=6.99 A=48.8601 P=27.96 m=1
C$123 \$45 VGND cap_cmim w=6.99 l=6.99 A=48.8601 P=27.96 m=1
C$124 Vout VGND cap_cmim w=6.99 l=6.99 A=48.8601 P=27.96 m=1
C$125 \$40 VGND cap_cmim w=6.99 l=6.99 A=48.8601 P=27.96 m=1
C$126 \$51 VGND cap_cmim w=6.99 l=6.99 A=48.8601 P=27.96 m=1
C$127 \$44 VGND cap_cmim w=6.99 l=6.99 A=48.8601 P=27.96 m=1
M$128 \$127 \$51 \$142 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$129 \$142 \$51 \$127 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
M$130 \$142 \$51 \$152 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.11
+ PS=0.945 PD=0.94
M$131 \$152 \$51 \$142 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.11 PS=0.94
+ PD=0.94
M$132 \$142 \$51 \$152 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
M$133 \$142 \$51 \$152 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.17
+ PS=0.945 PD=1.68
M$134 \$130 \$142 \$143 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$135 \$143 \$142 \$130 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
M$136 \$143 \$142 \$153 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.11
+ PS=0.945 PD=0.94
M$137 \$153 \$142 \$143 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.11 PS=0.94
+ PD=0.94
M$138 \$143 \$142 \$153 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
M$139 \$143 \$142 \$153 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.17
+ PS=0.945 PD=1.68
M$140 \$136 \$143 \$144 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$141 \$144 \$143 \$136 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
M$142 \$144 \$143 \$154 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.11
+ PS=0.945 PD=0.94
M$143 \$154 \$143 \$144 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.11 PS=0.94
+ PD=0.94
M$144 \$144 \$143 \$154 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
M$145 \$144 \$143 \$154 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.17
+ PS=0.945 PD=1.68
M$146 \$124 \$144 \$145 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$147 \$145 \$144 \$124 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
M$148 \$145 \$144 \$155 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.11
+ PS=0.945 PD=0.94
M$149 \$155 \$144 \$145 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.11 PS=0.94
+ PD=0.94
M$150 \$145 \$144 \$155 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
M$151 \$145 \$144 \$155 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.17
+ PS=0.945 PD=1.68
M$152 \$125 \$145 \$45 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.17 AD=0.11 PS=1.68
+ PD=0.94
M$153 \$45 \$145 \$125 VGND sg13_lv_nmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
M$154 \$45 \$145 \$156 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.11
+ PS=0.945 PD=0.94
M$155 \$156 \$145 \$45 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.11 PS=0.94
+ PD=0.94
M$156 \$45 \$145 \$156 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.11 AD=0.17 PS=0.94
+ PD=1.68
M$157 \$45 \$145 \$156 VPWR sg13_lv_pmos L=0.13 W=0.5 AS=0.1106 AD=0.17
+ PS=0.945 PD=1.68
.ENDS 11Stage_vco_new
