* Extracted by KLayout with SG13G2 LVS runset on : 12/08/2025 13:07

.SUBCKT pll_3bitDiv
X$1 1 1 20 2 16 18 10 10 Bias_gen
X$33602 1 2 3 10 5 6 12 7 3bit_freq_divider
X$35351 1 2 3 10 4 8 9 13 3bit_freq_divider
X$45101 10 1 20 2 sg13g2_inv_1
X$45828 1 10 11 12 17 14 PFD
X$48295 1 10 3 15 vco_wob
X$49096 17 11 18 16 10 19 1 charge_pump
X$49597 1 15 19 loop_filter
.ENDS pll_3bitDiv

.SUBCKT PFD 1 2 3 6 11 14
M$1 5 6 7 1 sg13_lv_nmos L=0.15u W=0.84u AS=0.2226p AD=0.2226p PS=2.32u PD=2.32u
M$3 10 14 12 1 sg13_lv_nmos L=0.15u W=0.84u AS=0.2226p AD=0.2226p PS=2.32u
+ PD=2.32u
M$5 1 13 11 1 sg13_lv_nmos L=0.15u W=0.48u AS=0.1632p AD=0.1632p PS=1.64u
+ PD=1.64u
M$6 1 4 3 1 sg13_lv_nmos L=0.15u W=0.48u AS=0.1632p AD=0.1632p PS=1.64u PD=1.64u
M$7 8 6 1 1 sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p PS=1.4u PD=1.4u
M$8 1 10 13 1 sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p PS=1.4u PD=1.4u
M$9 1 5 4 1 sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p PS=1.4u PD=1.4u
M$10 9 14 1 1 sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p PS=1.4u PD=1.4u
M$11 2 13 11 2 sg13_lv_pmos L=0.15u W=0.96u AS=0.2304p AD=0.2304p PS=2.72u
+ PD=2.72u
M$14 2 4 3 2 sg13_lv_pmos L=0.15u W=0.96u AS=0.2304p AD=0.2304p PS=2.72u
+ PD=2.72u
M$17 13 10 2 2 sg13_lv_pmos L=0.15u W=0.72u AS=0.1908p AD=0.1908p PS=2.14u
+ PD=2.14u
M$19 2 5 4 2 sg13_lv_pmos L=0.15u W=0.72u AS=0.1908p AD=0.1908p PS=2.14u
+ PD=2.14u
M$21 8 14 12 1 sg13_lv_nmos L=0.15u W=1.8u AS=0.396p AD=0.396p PS=4.36u PD=4.36u
M$26 9 6 7 1 sg13_lv_nmos L=0.15u W=1.8u AS=0.396p AD=0.396p PS=4.36u PD=4.36u
M$31 12 14 2 2 sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p AD=0.1696p PS=2.02u
+ PD=2.02u
M$33 7 6 2 2 sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p AD=0.1696p PS=2.02u
+ PD=2.02u
M$35 5 6 6 2 sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p AD=0.1696p PS=2.02u
+ PD=2.02u
M$37 10 14 14 2 sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p AD=0.1696p PS=2.02u
+ PD=2.02u
.ENDS PFD

.SUBCKT charge_pump 1 2 4 5 6 7 9
M$1 9 5 8 9 sg13_lv_nmos L=0.13u W=1.2u AS=0.408p AD=0.207p PS=3.08u PD=1.545u
M$2 8 2 7 9 sg13_lv_nmos L=0.13u W=1.2u AS=0.207p AD=0.408p PS=1.545u PD=3.08u
M$3 7 3 10 6 sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$4 10 4 6 6 sg13_lv_pmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$5 3 1 6 6 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u PD=1.28u
M$6 9 1 3 9 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u PD=1.34u
.ENDS charge_pump

.SUBCKT loop_filter 1 2 4
M$1 1 4 1 1 sg13_lv_nmos L=0.65u W=45u AS=9p AD=9p PS=60u PD=60u
R$31 4 2 rhigh w=0.6u l=0.96u ps=0 b=0 m=1
R$32 3 4 rhigh w=0.5u l=0.96u ps=0 b=0 m=1
M$33 1 2 1 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.201p AD=0.201p PS=2.68u PD=2.68u
M$35 1 3 1 1 sg13_lv_nmos L=0.65u W=15u AS=3p AD=3p PS=28u PD=28u
.ENDS loop_filter

.SUBCKT Bias_gen 1 2 4 5 6 9 10 13
R$1 11 13 rhigh w=1u l=12u ps=0 b=0 m=1
R$2 3 2 rhigh w=1u l=12u ps=0 b=0 m=1
M$3 7 6 2 1 sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$4 9 6 3 1 sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$5 6 6 2 1 sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$6 9 7 8 1 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
M$7 6 4 2 1 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
M$8 8 5 2 1 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
M$9 6 9 11 10 sg13_lv_pmos L=1u W=4u AS=1.06p AD=1.06p PS=7.06u PD=7.06u
M$11 13 9 9 10 sg13_lv_pmos L=1u W=2u AS=0.68p AD=0.68p PS=4.68u PD=4.68u
M$12 13 12 12 10 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
M$13 13 5 9 10 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
M$14 12 7 7 10 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
M$15 13 5 7 10 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
.ENDS Bias_gen

.SUBCKT vco_wob 1 2 12 23
M$1 18 14 13 1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u PD=2.62u
M$3 1 23 31 1 sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p PS=2.02u PD=2.02u
M$5 1 23 32 1 sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p PS=2.02u PD=2.02u
M$7 21 9 15 1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u PD=2.62u
M$9 19 11 14 1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u PD=2.62u
M$11 1 23 19 1 sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p PS=2.02u PD=2.02u
M$13 1 23 25 1 sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p PS=2.02u PD=2.02u
M$15 22 12 9 1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u PD=2.62u
M$17 1 23 10 1 sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p PS=2.02u PD=2.02u
M$19 20 15 11 1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u PD=2.62u
M$21 1 23 20 1 sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p PS=2.02u PD=2.02u
M$23 1 23 24 1 sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p PS=2.02u PD=2.02u
M$25 1 23 30 1 sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p PS=2.02u PD=2.02u
M$27 1 23 22 1 sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p PS=2.02u PD=2.02u
M$29 1 23 17 1 sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p PS=2.02u PD=2.02u
M$31 1 23 21 1 sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p PS=2.02u PD=2.02u
M$33 17 13 16 1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u PD=2.62u
M$35 1 23 18 1 sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p PS=2.02u PD=2.02u
M$37 3 10 2 2 sg13_lv_pmos L=0.13u W=0.8u AS=0.2825p AD=0.281p PS=3.57u PD=3.56u
M$41 4 10 2 2 sg13_lv_pmos L=0.13u W=0.8u AS=0.2825p AD=0.281p PS=3.57u PD=3.56u
M$45 11 15 5 2 sg13_lv_pmos L=0.13u W=2u AS=0.5012p AD=0.5p PS=4.51u PD=4.5u
M$49 6 10 2 2 sg13_lv_pmos L=0.13u W=0.8u AS=0.2825p AD=0.281p PS=3.57u PD=3.56u
M$53 8 10 2 2 sg13_lv_pmos L=0.13u W=0.8u AS=0.2825p AD=0.281p PS=3.57u PD=3.56u
M$57 7 10 2 2 sg13_lv_pmos L=0.13u W=0.8u AS=0.2825p AD=0.281p PS=3.57u PD=3.56u
M$61 16 13 3 2 sg13_lv_pmos L=0.13u W=2u AS=0.5012p AD=0.5p PS=4.51u PD=4.5u
M$65 5 10 2 2 sg13_lv_pmos L=0.13u W=0.8u AS=0.2825p AD=0.281p PS=3.57u PD=3.56u
M$69 2 10 10 2 sg13_lv_pmos L=0.13u W=0.8u AS=0.28175p AD=0.28175p PS=3.565u
+ PD=3.565u
M$73 34 10 2 2 sg13_lv_pmos L=0.13u W=0.8u AS=0.2375p AD=0.326p PS=2.97u
+ PD=4.16u
M$77 35 10 2 2 sg13_lv_pmos L=0.13u W=0.8u AS=0.2375p AD=0.326p PS=2.97u
+ PD=4.16u
M$81 14 11 4 2 sg13_lv_pmos L=0.13u W=2u AS=0.5012p AD=0.5p PS=4.51u PD=4.5u
M$85 9 12 7 2 sg13_lv_pmos L=0.13u W=2u AS=0.5012p AD=0.5p PS=4.51u PD=4.5u
M$89 15 9 6 2 sg13_lv_pmos L=0.13u W=2u AS=0.5012p AD=0.5p PS=4.51u PD=4.5u
M$93 33 10 2 2 sg13_lv_pmos L=0.13u W=0.8u AS=0.2375p AD=0.326p PS=2.97u
+ PD=4.16u
M$97 13 14 8 2 sg13_lv_pmos L=0.13u W=2u AS=0.5012p AD=0.5p PS=4.51u PD=4.5u
M$101 36 10 2 2 sg13_lv_pmos L=0.13u W=0.8u AS=0.2375p AD=0.326p PS=2.97u
+ PD=4.16u
M$105 37 10 2 2 sg13_lv_pmos L=0.13u W=0.8u AS=0.2375p AD=0.326p PS=2.97u
+ PD=4.16u
C$109 14 1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$110 27 1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$111 29 1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$112 26 1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$113 15 1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$114 11 1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$115 9 1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$116 13 1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$117 28 1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$118 12 1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$119 16 1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
M$120 30 16 26 1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u PD=2.62u
M$122 26 16 33 2 sg13_lv_pmos L=0.13u W=2u AS=0.4412p AD=0.56p PS=3.77u PD=5.24u
M$126 31 26 27 1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u PD=2.62u
M$128 27 26 34 2 sg13_lv_pmos L=0.13u W=2u AS=0.4412p AD=0.56p PS=3.77u PD=5.24u
M$132 32 27 28 1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u PD=2.62u
M$134 28 27 35 2 sg13_lv_pmos L=0.13u W=2u AS=0.4412p AD=0.56p PS=3.77u PD=5.24u
M$138 24 28 29 1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u PD=2.62u
M$140 29 28 36 2 sg13_lv_pmos L=0.13u W=2u AS=0.4412p AD=0.56p PS=3.77u PD=5.24u
M$144 25 29 12 1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u PD=2.62u
M$146 12 29 37 2 sg13_lv_pmos L=0.13u W=2u AS=0.4412p AD=0.56p PS=3.77u PD=5.24u
.ENDS vco_wob

.SUBCKT 3bit_freq_divider 1 2 3 5 10 12 15 17
X$1 13 5 1 sg13g2_tiehi
X$2 6 11 11 15 1 13 5 dff_nclk
X$3 5 1 8 9 7 6 sg13g2_or3_1
X$4 16 14 4 12 7 6 1 5 freq_div_cell
X$5 18 16 4 17 8 6 1 5 freq_div_cell
X$6 18 5 1 sg13g2_tiehi
X$7 14 19 4 10 9 6 1 5 freq_div_cell
X$8 5 1 4 3 2 sg13g2_nand2_1
.ENDS 3bit_freq_divider

.SUBCKT sg13g2_nand2_1 1 2 3 4 5
M$1 2 5 6 2 sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.0666p PS=2.16u PD=0.92u
M$2 6 4 3 2 sg13_lv_nmos L=0.13u W=0.74u AS=0.0666p AD=0.2516p PS=0.92u PD=2.16u
M$3 1 5 3 1 sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.2128p PS=2.92u PD=1.5u
M$4 3 4 1 1 sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.3808p PS=1.5u PD=2.92u
.ENDS sg13g2_nand2_1

.SUBCKT sg13g2_or3_1 1 2 3 4 5 7
M$1 6 3 2 2 sg13_lv_nmos L=0.13u W=0.55u AS=0.187p AD=0.1045p PS=1.78u PD=0.93u
M$2 2 5 6 2 sg13_lv_nmos L=0.13u W=0.55u AS=0.1045p AD=0.198p PS=0.93u PD=1.27u
M$3 6 4 2 2 sg13_lv_nmos L=0.13u W=0.55u AS=0.198p AD=0.13395p PS=1.27u PD=1.12u
M$4 2 6 7 2 sg13_lv_nmos L=0.13u W=0.74u AS=0.13395p AD=0.2516p PS=1.12u
+ PD=2.16u
M$5 6 3 9 1 sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.1275p PS=2.68u PD=1.255u
M$6 9 5 8 1 sg13_lv_pmos L=0.13u W=1u AS=0.1275p AD=0.22p PS=1.255u PD=1.44u
M$7 8 4 1 1 sg13_lv_pmos L=0.13u W=1u AS=0.22p AD=0.3822p PS=1.44u PD=1.84u
M$8 1 6 7 1 sg13_lv_pmos L=0.13u W=1.12u AS=0.3822p AD=0.3808p PS=1.84u PD=2.92u
.ENDS sg13g2_or3_1

.SUBCKT sg13g2_tiehi 2 5 6
M$1 6 4 4 6 sg13_lv_nmos L=0.13u W=0.3u AS=0.2307p AD=0.102p PS=1.615u PD=1.28u
M$2 6 3 1 6 sg13_lv_nmos L=0.13u W=0.795u AS=0.2307p AD=0.274275p PS=1.615u
+ PD=2.28u
M$3 3 4 5 5 sg13_lv_pmos L=0.13u W=0.66u AS=0.2442p AD=0.4657125p PS=2.06u
+ PD=2.54u
M$4 5 1 2 5 sg13_lv_pmos L=0.13u W=1.155u AS=0.4657125p AD=0.3927p PS=2.54u
+ PD=2.99u
.ENDS sg13g2_tiehi

.SUBCKT freq_div_cell 1 2 3 4 5 7 9 10
X$1 1 6 8 2 9 10 half_add
X$2 3 8 11 6 9 7 10 dff_nclk
X$3 9 5 10 6 4 sg13g2_xor2_1
.ENDS freq_div_cell

.SUBCKT dff_nclk 1 2 3 4 6 7 8
X$1 8 6 1 5 sg13g2_inv_1
X$2 6 7 3 4 2 5 8 sg13g2_dfrbp_1
.ENDS dff_nclk

.SUBCKT half_add 1 2 3 4 5 6
X$1 5 3 6 1 2 sg13g2_xor2_1
X$2 6 5 4 1 2 sg13g2_and2_1
.ENDS half_add

.SUBCKT sg13g2_dfrbp_1 1 2 7 9 10 12 20
M$1 5 11 19 1 sg13_lv_nmos L=0.13u W=0.42u AS=0.2017p AD=0.0546p PS=1.48u
+ PD=0.68u
M$2 19 6 1 1 sg13_lv_nmos L=0.13u W=0.42u AS=0.0546p AD=0.0903p PS=0.68u
+ PD=0.85u
M$3 1 2 18 1 sg13_lv_nmos L=0.13u W=0.42u AS=0.0903p AD=0.04725p PS=0.85u
+ PD=0.645u
M$4 18 5 6 1 sg13_lv_nmos L=0.13u W=0.42u AS=0.04725p AD=0.1428p PS=0.645u
+ PD=1.52u
M$5 1 13 14 1 sg13_lv_nmos L=0.13u W=0.64u AS=0.1825p AD=0.193975p PS=1.325u
+ PD=1.29u
M$6 14 3 5 1 sg13_lv_nmos L=0.13u W=0.64u AS=0.193975p AD=0.2017p PS=1.29u
+ PD=1.48u
M$7 4 11 13 1 sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p PS=1.52u
+ PD=0.8u
M$8 13 3 16 1 sg13_lv_nmos L=0.13u W=0.42u AS=0.0798p AD=0.0546p PS=0.8u
+ PD=0.68u
M$9 16 14 17 1 sg13_lv_nmos L=0.13u W=0.42u AS=0.0546p AD=0.0483p PS=0.68u
+ PD=0.65u
M$10 1 2 17 1 sg13_lv_nmos L=0.13u W=0.42u AS=0.1825p AD=0.0483p PS=1.325u
+ PD=0.65u
M$11 8 5 1 1 sg13_lv_nmos L=0.13u W=0.55u AS=0.187p AD=0.14505p PS=1.78u
+ PD=1.15u
M$12 1 8 9 1 sg13_lv_nmos L=0.13u W=0.74u AS=0.14505p AD=0.2516p PS=1.15u
+ PD=2.16u
M$13 1 5 7 1 sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.2775p PS=2.16u
+ PD=2.23u
M$14 1 12 11 1 sg13_lv_nmos L=0.13u W=0.74u AS=0.1544p AD=0.2516p PS=1.235u
+ PD=2.16u
M$15 1 11 3 1 sg13_lv_nmos L=0.13u W=0.74u AS=0.1544p AD=0.2516p PS=1.235u
+ PD=2.16u
M$16 4 10 15 1 sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.0504p PS=1.52u
+ PD=0.66u
M$17 15 2 1 1 sg13_lv_nmos L=0.13u W=0.42u AS=0.0504p AD=0.1428p PS=0.66u
+ PD=1.52u
M$18 11 12 20 20 sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.19p PS=2.68u PD=1.38u
M$19 20 11 3 20 sg13_lv_pmos L=0.13u W=1u AS=0.19p AD=0.34p PS=1.38u PD=2.68u
M$20 20 10 4 20 sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p PS=1.52u
+ PD=0.8u
M$21 4 2 20 20 sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.1428p PS=0.8u
+ PD=1.52u
M$22 20 5 8 20 sg13_lv_pmos L=0.13u W=0.84u AS=0.2016p AD=0.2856p PS=1.5u
+ PD=2.36u
M$23 20 8 9 20 sg13_lv_pmos L=0.13u W=1.12u AS=0.2016p AD=0.3808p PS=1.5u
+ PD=2.92u
M$24 20 13 14 20 sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.19p PS=2.68u PD=1.38u
M$25 14 11 5 20 sg13_lv_pmos L=0.13u W=1u AS=0.19p AD=0.17695p PS=1.38u PD=1.56u
M$26 5 3 22 20 sg13_lv_pmos L=0.13u W=0.42u AS=0.17695p AD=0.04305p PS=1.56u
+ PD=0.625u
M$27 22 6 20 20 sg13_lv_pmos L=0.13u W=0.42u AS=0.04305p AD=0.0798p PS=0.625u
+ PD=0.8u
M$28 20 2 6 20 sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.0798p PS=0.8u
+ PD=0.8u
M$29 20 5 6 20 sg13_lv_pmos L=0.13u W=0.42u AS=0.2163p AD=0.0798p PS=1.55u
+ PD=0.8u
M$30 20 5 7 20 sg13_lv_pmos L=0.13u W=1.12u AS=0.2163p AD=0.7616p PS=1.55u
+ PD=3.6u
M$31 4 3 13 20 sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p PS=1.52u
+ PD=0.8u
M$32 13 11 21 20 sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.05145p PS=0.8u
+ PD=0.665u
M$33 21 14 20 20 sg13_lv_pmos L=0.13u W=0.42u AS=0.05145p AD=0.11785p PS=0.665u
+ PD=1.025u
M$34 20 2 13 20 sg13_lv_pmos L=0.13u W=0.42u AS=0.11785p AD=0.1533p PS=1.025u
+ PD=1.57u
.ENDS sg13g2_dfrbp_1

.SUBCKT sg13g2_inv_1 1 2 3 4
M$1 2 3 4 2 sg13_lv_nmos L=0.13u W=0.74u AS=0.259p AD=0.259p PS=2.18u PD=2.18u
M$2 1 3 4 1 sg13_lv_pmos L=0.13u W=1.12u AS=0.392p AD=0.392p PS=2.94u PD=2.94u
.ENDS sg13g2_inv_1

.SUBCKT sg13g2_and2_1 1 2 3 4 5
M$1 6 4 7 2 sg13_lv_nmos L=0.13u W=0.64u AS=0.2176p AD=0.1216p PS=1.96u PD=1.02u
M$2 2 5 7 2 sg13_lv_nmos L=0.13u W=0.64u AS=0.1331p AD=0.1216p PS=1.12u PD=1.02u
M$3 2 6 3 2 sg13_lv_nmos L=0.13u W=0.74u AS=0.1331p AD=0.2516p PS=1.12u PD=2.16u
M$4 1 4 6 1 sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p AD=0.1596p PS=2.36u PD=1.22u
M$5 1 5 6 1 sg13_lv_pmos L=0.13u W=0.84u AS=0.1918p AD=0.1596p PS=1.5u PD=1.22u
M$6 1 6 3 1 sg13_lv_pmos L=0.13u W=1.12u AS=0.1918p AD=0.3808p PS=1.5u PD=2.92u
.ENDS sg13g2_and2_1

.SUBCKT sg13g2_xor2_1 2 4 5 6 7
M$1 2 6 1 2 sg13_lv_nmos L=0.13u W=0.55u AS=0.374p AD=0.174625p PS=2.46u
+ PD=1.185u
M$2 2 7 1 2 sg13_lv_nmos L=0.13u W=0.55u AS=0.15245p AD=0.174625p PS=1.17u
+ PD=1.185u
M$3 2 6 8 2 sg13_lv_nmos L=0.13u W=0.74u AS=0.15245p AD=0.0888p PS=1.17u
+ PD=0.98u
M$4 8 7 4 2 sg13_lv_nmos L=0.13u W=0.74u AS=0.0888p AD=0.1628p PS=0.98u PD=1.18u
M$5 4 1 2 2 sg13_lv_nmos L=0.13u W=0.74u AS=0.1628p AD=0.3108p PS=1.18u PD=2.32u
M$6 3 6 5 5 sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.2128p PS=2.92u PD=1.5u
M$7 5 7 3 5 sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.2128p PS=1.5u PD=1.5u
M$8 3 1 4 5 sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.3808p PS=1.5u PD=2.92u
M$9 5 6 9 5 sg13_lv_pmos L=0.13u W=1u AS=0.36p AD=0.1225p PS=2.72u PD=1.245u
M$10 9 7 1 5 sg13_lv_pmos L=0.13u W=1u AS=0.1225p AD=0.34p PS=1.245u PD=2.68u
.ENDS sg13g2_xor2_1
