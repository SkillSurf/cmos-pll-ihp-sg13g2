* Extracted by KLayout with SG13G2 LVS runset on : 11/06/2025 12:36

.SUBCKT t2_vco_new
M$1 1 3 4 1 sg13_lv_nmos L=0.13u W=1u AS=0.295p AD=0.295p PS=3.56u PD=3.56u
M$5 1 3 5 1 sg13_lv_nmos L=0.13u W=1u AS=0.295p AD=0.295p PS=3.56u PD=3.56u
M$9 1 3 6 1 sg13_lv_nmos L=0.13u W=1u AS=0.295p AD=0.295p PS=3.56u PD=3.56u
M$13 1 3 7 1 sg13_lv_nmos L=0.13u W=1u AS=0.295p AD=0.295p PS=3.56u PD=3.56u
M$17 1 3 8 1 sg13_lv_nmos L=0.13u W=1u AS=0.295p AD=0.295p PS=3.56u PD=3.56u
M$21 1 3 9 1 sg13_lv_nmos L=0.13u W=1u AS=0.295p AD=0.295p PS=3.56u PD=3.56u
M$25 5 2 10 1 sg13_lv_nmos L=0.13u W=0.5u AS=0.17p AD=0.17p PS=2.08u PD=2.08u
M$27 6 10 11 1 sg13_lv_nmos L=0.13u W=0.5u AS=0.17p AD=0.17p PS=2.08u PD=2.08u
M$29 7 11 12 1 sg13_lv_nmos L=0.13u W=0.5u AS=0.17p AD=0.17p PS=2.08u PD=2.08u
M$31 8 12 13 1 sg13_lv_nmos L=0.13u W=0.5u AS=0.17p AD=0.17p PS=2.08u PD=2.08u
M$33 9 13 14 1 sg13_lv_nmos L=0.13u W=0.5u AS=0.17p AD=0.17p PS=2.08u PD=2.08u
M$35 1 14 2 1 sg13_lv_nmos L=0.13u W=0.5u AS=0.17p AD=0.17p PS=2.08u PD=2.08u
M$37 10 2 4 16 sg13_lv_pmos L=0.13u W=1u AS=0.2515p AD=0.34p PS=2.97u PD=4.16u
M$41 11 10 4 18 sg13_lv_pmos L=0.13u W=1u AS=0.2515p AD=0.34p PS=2.97u PD=4.16u
M$45 12 11 4 19 sg13_lv_pmos L=0.13u W=1u AS=0.2515p AD=0.34p PS=2.97u PD=4.16u
M$49 13 12 4 20 sg13_lv_pmos L=0.13u W=1u AS=0.2515p AD=0.34p PS=2.97u PD=4.16u
M$53 14 13 4 17 sg13_lv_pmos L=0.13u W=1u AS=0.2515p AD=0.34p PS=2.97u PD=4.16u
M$57 2 14 4 15 sg13_lv_pmos L=0.13u W=1u AS=0.2515p AD=0.34p PS=2.97u PD=4.16u
.ENDS t2_vco_new
