** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_inverter_tb_dc.sch
**.subckt t2_inverter_tb_dc Vout
*.opin Vout
Vin Vin GND 0
Vdd Vdd GND 1.2
x1 Vdd Vin Vout GND t2_inverter
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt




.param temp=27
.control
dc Vin 0 1.2 0.1
.save all
plot v(Vin) v(Vout)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/IHP/Inverter/t2_inverter.sym # of pins=4
** sym_path: /foss/designs/IHP/Inverter/t2_inverter.sym
** sch_path: /foss/designs/IHP/Inverter/t2_inverter.sch
.subckt t2_inverter VP A Y VN
*.iopin VP
*.iopin VN
*.ipin A
*.opin Y
XM2 Y A VP VP sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
XM1 Y A VN VN sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
