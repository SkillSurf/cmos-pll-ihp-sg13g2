* Extracted by KLayout with SG13G2 LVS runset on : 13/06/2025 00:18

.SUBCKT t2_bais
M$1 3 3 4 1 sg13_lv_nmos L=1u W=0.2u AS=0.104p AD=0.059p PS=1.34u PD=0.74u
M$2 4 3 3 1 sg13_lv_nmos L=1u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$3 3 3 4 1 sg13_lv_nmos L=1u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$4 4 3 3 1 sg13_lv_nmos L=1u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$5 3 3 4 1 sg13_lv_nmos L=1u W=0.2u AS=0.059p AD=0.104p PS=0.74u PD=1.34u
M$6 3 3 3 1 sg13_lv_nmos L=1u W=0.2u AS=0.104p AD=0.059p PS=1.34u PD=0.74u
M$7 3 3 3 1 sg13_lv_nmos L=1u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$8 3 3 3 1 sg13_lv_nmos L=1u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$9 3 3 3 1 sg13_lv_nmos L=1u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$10 3 3 3 1 sg13_lv_nmos L=1u W=0.2u AS=0.059p AD=0.104p PS=0.74u PD=1.34u
M$11 4 3 6 1 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.095p PS=1.68u PD=0.88u
M$12 6 5 7 1 sg13_lv_nmos L=0.15u W=0.5u AS=0.095p AD=0.17p PS=0.88u PD=1.68u
M$13 3 2 3 1 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
M$14 3 3 11 8 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.095p PS=1.68u PD=0.88u
M$15 11 11 10 8 sg13_lv_pmos L=0.15u W=0.5u AS=0.095p AD=0.17p PS=0.88u PD=1.68u
M$16 3 5 10 8 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
M$17 3 5 10 8 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
M$18 10 3 3 8 sg13_lv_pmos L=1u W=0.2u AS=0.104p AD=0.059p PS=1.34u PD=0.74u
M$19 3 3 10 8 sg13_lv_pmos L=1u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$20 10 3 3 8 sg13_lv_pmos L=1u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$21 3 3 10 8 sg13_lv_pmos L=1u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$22 10 3 3 8 sg13_lv_pmos L=1u W=0.2u AS=0.059p AD=0.104p PS=0.74u PD=1.34u
M$23 9 3 3 8 sg13_lv_pmos L=1u W=0.2u AS=0.104p AD=0.059p PS=1.34u PD=0.74u
M$24 3 3 9 8 sg13_lv_pmos L=1u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$25 9 3 3 8 sg13_lv_pmos L=1u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$26 3 3 9 8 sg13_lv_pmos L=1u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$27 9 3 3 8 sg13_lv_pmos L=1u W=0.2u AS=0.059p AD=0.104p PS=0.74u PD=1.34u
R$28 9 10 rhigh w=0.5u l=0.5u ps=0 b=0 m=1
.ENDS t2_bais
