** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_vco_new.sch
.subckt t2_vco_new VPWR VGND vctl Vout
*.PININFO VPWR:B VGND:B vctl:I Vout:O
M1 mirror_pg mirror_pg VPWR VPWR sg13_lv_pmos w=2u l=0.13u ng=1 m=1
M2 net1 mirror_pg VPWR VPWR sg13_lv_pmos w=2u l=0.13u ng=1 m=1
M3 net2 mirror_pg VPWR VPWR sg13_lv_pmos w=2u l=0.13u ng=1 m=1
M4 net3 mirror_pg VPWR VPWR sg13_lv_pmos w=2u l=0.13u ng=1 m=1
M5 mirror_pg vctl VGND VGND sg13_lv_nmos w=1u l=0.13u ng=1 m=1
M6 net9 vctl VGND VGND sg13_lv_nmos w=1u l=0.13u ng=1 m=1
M7 net8 vctl VGND VGND sg13_lv_nmos w=1u l=0.13u ng=1 m=1
M8 net7 vctl VGND VGND sg13_lv_nmos w=1u l=0.13u ng=1 m=1
C1 feedback VGND 10f m=1
C2 Vout VGND 20f m=1
M9 net13 mirror_pg VPWR VPWR sg13_lv_pmos w=2u l=0.13u ng=1 m=1
M10 net12 mirror_pg VPWR VPWR sg13_lv_pmos w=2u l=0.13u ng=1 m=1
M11 net10 vctl VGND VGND sg13_lv_nmos w=1u l=0.13u ng=1 m=1
M12 net11 vctl VGND VGND sg13_lv_nmos w=1u l=0.13u ng=1 m=1
x7 net1 VPWR feedback net4 VGND net9 t2_vco_inverter
x1 net2 VPWR net4 net5 VGND net8 t2_vco_inverter
x2 net3 VPWR net5 net6 VGND net7 t2_vco_inverter
x3 net13 VPWR net6 net14 VGND net10 t2_vco_inverter
x4 net12 VPWR net14 feedback VGND net11 t2_vco_inverter
x5 VPWR VPWR feedback Vout VGND VGND t2_vco_inverter
.ends

* expanding   symbol:  t2_vco_inverter.sym # of pins=6
** sym_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_vco_inverter.sym
** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_vco_inverter.sch
.subckt t2_vco_inverter VPWR VPB A Y VNB VGND
*.PININFO VPWR:B VGND:B A:I Y:O VPB:B VNB:B
M2 Y A VPWR VPB sg13_lv_pmos w=1u l=0.13u ng=1 m=1
M1 Y A VGND VNB sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
.ends

