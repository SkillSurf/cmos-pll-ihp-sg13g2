* Extracted by KLayout with SG13G2 LVS runset on : 10/06/2025 18:05

.SUBCKT t2_inverter
M$1 1 4 3 1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u PD=1.34u
M$2 2 4 3 2 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u PD=1.28u
.ENDS t2_inverter
