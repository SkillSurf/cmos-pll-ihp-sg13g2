* Extracted by KLayout with SG13G2 LVS runset on : 13/07/2025 07:28

.SUBCKT PFD VDD VSS DOWN VCO_CLK UP Ref_CLK
M$1 \$5 VCO_CLK \$7 VSS sg13_lv_nmos L=0.15u W=0.84u AS=0.2226p AD=0.2226p
+ PS=2.32u PD=2.32u
M$3 \$10 Ref_CLK \$12 VSS sg13_lv_nmos L=0.15u W=0.84u AS=0.2226p AD=0.2226p
+ PS=2.32u PD=2.32u
M$5 VSS \$13 UP VSS sg13_lv_nmos L=0.15u W=0.48u AS=0.1632p AD=0.1632p PS=1.64u
+ PD=1.64u
M$6 VSS \$4 DOWN VSS sg13_lv_nmos L=0.15u W=0.48u AS=0.1632p AD=0.1632p
+ PS=1.64u PD=1.64u
M$7 \$8 VCO_CLK VSS VSS sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p
+ PS=1.4u PD=1.4u
M$8 VSS \$10 \$13 VSS sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p
+ PS=1.4u PD=1.4u
M$9 VSS \$5 \$4 VSS sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p PS=1.4u
+ PD=1.4u
M$10 \$9 Ref_CLK VSS VSS sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p
+ PS=1.4u PD=1.4u
M$11 VDD \$13 UP VDD sg13_lv_pmos L=0.15u W=0.96u AS=0.2304p AD=0.2304p
+ PS=2.72u PD=2.72u
M$14 VDD \$4 DOWN VDD sg13_lv_pmos L=0.15u W=0.96u AS=0.2304p AD=0.2304p
+ PS=2.72u PD=2.72u
M$17 \$13 \$10 VDD VDD sg13_lv_pmos L=0.15u W=0.72u AS=0.1908p AD=0.1908p
+ PS=2.14u PD=2.14u
M$19 VDD \$5 \$4 VDD sg13_lv_pmos L=0.15u W=0.72u AS=0.1908p AD=0.1908p
+ PS=2.14u PD=2.14u
M$21 \$8 Ref_CLK \$12 VSS sg13_lv_nmos L=0.15u W=1.8u AS=0.396p AD=0.396p
+ PS=4.36u PD=4.36u
M$26 \$9 VCO_CLK \$7 VSS sg13_lv_nmos L=0.15u W=1.8u AS=0.396p AD=0.396p
+ PS=4.36u PD=4.36u
M$31 \$12 Ref_CLK VDD VDD sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p AD=0.1696p
+ PS=2.02u PD=2.02u
M$33 \$7 VCO_CLK VDD VDD sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p AD=0.1696p
+ PS=2.02u PD=2.02u
M$35 \$5 VCO_CLK VCO_CLK VDD sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p AD=0.1696p
+ PS=2.02u PD=2.02u
M$37 \$10 Ref_CLK Ref_CLK VDD sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p
+ AD=0.1696p PS=2.02u PD=2.02u
.ENDS PFD
