* Extracted by KLayout with SG13G2 LVS runset on : 10/06/2025 18:01

.SUBCKT t2_nand3
M$1 3 2 4 1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u PD=0.74u
M$2 4 5 6 1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p PS=0.74u PD=0.74u
M$3 6 7 1 1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u PD=1.34u
M$4 8 2 3 8 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$5 3 5 8 8 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.057p PS=0.68u PD=0.68u
M$6 8 7 3 8 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u PD=1.28u
.ENDS t2_nand3
