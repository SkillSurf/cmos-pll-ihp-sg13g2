* Extracted by KLayout with SG13G2 LVS runset on : 13/06/2025 12:35

.SUBCKT t2_charge_pump.gds
X$1 5 9 5 1 nmos$3
X$2 9 7 5 2 nmos$3
X$3 8 5 3 t2_inverter
X$4 7 10 3 6 5 pmos$2
X$5 10 8 4 6 5 pmos
M$1 5 1 9 5 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u PD=0.74u
M$2 9 2 7 5 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u PD=1.34u
M$3 7 3 10 6 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.05625p PS=1.28u PD=0.71u
M$4 10 4 8 6 sg13_lv_pmos L=0.13u W=0.15u AS=0.05625p AD=0.1005p PS=0.71u
+ PD=1.34u
.ENDS t2_charge_pump.gds

.SUBCKT pmos 1 2 3 4 5
.ENDS pmos

.SUBCKT pmos$2 1 2 3 4 5
.ENDS pmos$2

.SUBCKT nmos$3 1 2 3 4
.ENDS nmos$3

.SUBCKT t2_inverter 1 2 4
X$1 1 4 3 1 2 pmos$1
X$2 2 4 2 3 nmos
.ENDS t2_inverter

.SUBCKT pmos$1 1 2 3 4 5
M$1 1 3 2 4 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u PD=1.28u
.ENDS pmos$1

.SUBCKT nmos 1 2 3 4
M$1 1 4 2 3 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u PD=1.34u
.ENDS nmos
