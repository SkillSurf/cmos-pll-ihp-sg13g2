* Extracted by KLayout with SG13G2 LVS runset on : 11/06/2025 06:55

.SUBCKT t2_dff
X$1 2 4 10 1 12 t2_nand2
X$2 1 10 6 7 4 2 t2_nand3
X$3 2 1 9 7 t2_inverter
X$4 1 12 10 7 3 2 t2_nand3
X$5 1 11 8 6 3 2 t2_nand3
X$6 1 6 4 5 3 2 t2_nand3
X$7 2 10 8 1 11 t2_nand2
.ENDS t2_dff

.SUBCKT t2_inverter 1 2 3 4
M$1 1 3 4 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u PD=1.28u
M$2 2 3 4 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u PD=1.34u
.ENDS t2_inverter

.SUBCKT t2_nand3 1 2 3 4 5 8
M$1 3 2 6 1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u PD=0.74u
M$2 6 4 7 1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p PS=0.74u PD=0.74u
M$3 7 5 1 1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u PD=1.34u
M$4 8 2 3 8 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$5 3 4 8 8 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.057p PS=0.68u PD=0.68u
M$6 8 5 3 8 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u PD=1.28u
.ENDS t2_nand3

.SUBCKT t2_nand2 1 2 3 4 5
M$1 4 2 6 4 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u PD=0.74u
M$2 6 3 5 4 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u PD=1.34u
M$3 1 2 5 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$4 5 3 1 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u PD=1.28u
.ENDS t2_nand2
