** sch_path: /foss/designs/Team2/inverter/inverter.sch
**.subckt inverter VP A Y VN
*.iopin VN
*.iopin VP
*.ipin A
*.opin Y
XM1 Y A VP VP sg13_lv_pmos w=2u l=0.13u ng=1 m=1 rfmode=1
XM2 Y A VN VN sg13_lv_nmos w=1u l=0.13u ng=1 m=1 rfmode=1
**.ends
.end
