** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Combined_Design/design_data/xschem/2bit_freq_divider_pex_tb.sch

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.include ../../pex/2bit_freq_divider__2bit_freq_divider/magic_RC/2bit_freq_divider.pex.spice

**.subckt 2bit_freq_divider_pex_tb
Vs VDD GND 1.2
Vclk CLK_IN GND dc 0 ac 0 pulse(0, 1.2, 0, 100p, 100p, 6.25n, 12.5n)
* noconn CLK_OUT
Ven EN GND dc {EN}
Va0 A0 GND dc {A0}
Va1 A1 GND dc {A1}
x1 VDD GND A0 CLK_OUT CLK_IN EN A1 2bit_freq_divider
**** begin user architecture code


.meas tran tperiod_in TRIG v(clk_in) VAL=0.5 FALL=1 TARG v(clk_in) VAL=0.5 FALL=2
.meas tran freq_in PARAM = '1e-6/tperiod_in'

.meas tran tperiod_out TRIG v(clk_out) VAL=0.5 FALL=1 TARG v(clk_out) VAL=0.5 FALL=2
.meas tran freq_out PARAM = '1e-6/tperiod_out'

.meas tran tdelay TRIG v(clk_in) VAL=0.5 RISE=1 TARG v(clk_out) VAL=0.5 RISE=1




.param EN = 1.2

.param A0 = 1.2
.param A1 = 1.2




.param temp=27

.control
save all
tran 50p 150n

write tran_2bit_freq_divider_pex.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
