* Extracted by KLayout with SG13G2 LVS runset on : 10/06/2025 18:08

.SUBCKT t2_and2
M$1 4 3 5 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u PD=0.74u
M$2 5 8 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u PD=1.34u
M$3 6 4 7 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u PD=0.74u
M$4 7 4 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u PD=1.34u
M$5 1 3 4 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$6 4 8 1 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$7 1 4 6 1 sg13_lv_pmos L=0.13u W=0.6u AS=0.159p AD=0.159p PS=1.96u PD=1.96u
.ENDS t2_and2
