* Extracted by KLayout with SG13G2 LVS runset on : 13/06/2025 12:40

.SUBCKT t2_charge_pump
X$3 8 5 3 t2_inverter
M$1 5 1 10 5 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$2 10 2 7 5 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$3 7 3 9 6 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.05625p PS=1.28u PD=0.71u
M$4 9 4 8 6 sg13_lv_pmos L=0.13u W=0.15u AS=0.05625p AD=0.1005p PS=0.71u
+ PD=1.34u
.ENDS t2_charge_pump

.SUBCKT t2_inverter 1 2 4
M$1 1 3 4 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u PD=1.28u
M$2 2 3 4 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u PD=1.34u
.ENDS t2_inverter
