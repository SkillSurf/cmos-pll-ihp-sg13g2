* Extracted by KLayout with SG13G2 LVS runset on : 12/07/2025 14:50

.SUBCKT PFD
M$1 \$2 \$44 \$30 \$2 sg13_lv_nmos L=0.15u W=0.48u AS=0.1632p AD=0.1632p
+ PS=1.64u PD=1.64u
M$2 \$2 \$6 \$3 \$2 sg13_lv_nmos L=0.15u W=0.48u AS=0.1632p AD=0.1632p PS=1.64u
+ PD=1.64u
M$3 \$42 \$41 \$39 \$2 sg13_lv_nmos L=0.15u W=0.42u AS=0.1428p AD=0.0798p
+ PS=1.52u PD=0.8u
M$4 \$39 \$41 \$43 \$2 sg13_lv_nmos L=0.15u W=0.42u AS=0.0798p AD=0.1428p
+ PS=0.8u PD=1.52u
M$5 \$17 \$8 \$25 \$2 sg13_lv_nmos L=0.15u W=0.42u AS=0.1428p AD=0.0798p
+ PS=1.52u PD=0.8u
M$6 \$25 \$8 \$7 \$2 sg13_lv_nmos L=0.15u W=0.42u AS=0.0798p AD=0.1428p PS=0.8u
+ PD=1.52u
M$7 \$18 \$8 \$2 \$2 sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p PS=1.4u
+ PD=1.4u
M$8 \$2 \$43 \$44 \$2 sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p
+ PS=1.4u PD=1.4u
M$9 \$2 \$7 \$6 \$2 sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p PS=1.4u
+ PD=1.4u
M$10 \$19 \$41 \$2 \$2 sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p
+ PS=1.4u PD=1.4u
M$11 \$1 \$44 \$45 \$1 sg13_lv_pmos L=0.15u W=0.32u AS=0.1088p AD=0.0608p
+ PS=1.32u PD=0.7u
M$12 \$45 \$44 \$48 \$1 sg13_lv_pmos L=0.15u W=0.32u AS=0.0608p AD=0.0608p
+ PS=0.7u PD=0.7u
M$13 \$48 \$44 \$30 \$1 sg13_lv_pmos L=0.15u W=0.32u AS=0.0608p AD=0.1088p
+ PS=0.7u PD=1.32u
M$14 \$1 \$6 \$9 \$1 sg13_lv_pmos L=0.15u W=0.32u AS=0.1088p AD=0.0608p
+ PS=1.32u PD=0.7u
M$15 \$9 \$6 \$11 \$1 sg13_lv_pmos L=0.15u W=0.32u AS=0.0608p AD=0.0608p
+ PS=0.7u PD=0.7u
M$16 \$11 \$6 \$3 \$1 sg13_lv_pmos L=0.15u W=0.32u AS=0.0608p AD=0.1088p
+ PS=0.7u PD=1.32u
M$17 \$1 \$43 \$53 \$1 sg13_lv_pmos L=0.15u W=0.36u AS=0.1224p AD=0.0684p
+ PS=1.4u PD=0.74u
M$18 \$53 \$43 \$44 \$1 sg13_lv_pmos L=0.15u W=0.36u AS=0.0684p AD=0.1224p
+ PS=0.74u PD=1.4u
M$19 \$1 \$7 \$13 \$1 sg13_lv_pmos L=0.15u W=0.36u AS=0.1224p AD=0.0684p
+ PS=1.4u PD=0.74u
M$20 \$13 \$7 \$6 \$1 sg13_lv_pmos L=0.15u W=0.36u AS=0.0684p AD=0.1224p
+ PS=0.74u PD=1.4u
M$21 \$18 \$41 \$34 \$2 sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.0684p
+ PS=1.4u PD=0.74u
M$22 \$34 \$41 \$36 \$2 sg13_lv_nmos L=0.15u W=0.36u AS=0.0684p AD=0.0684p
+ PS=0.74u PD=0.74u
M$23 \$36 \$41 \$32 \$2 sg13_lv_nmos L=0.15u W=0.36u AS=0.0684p AD=0.0684p
+ PS=0.74u PD=0.74u
M$24 \$32 \$41 \$31 \$2 sg13_lv_nmos L=0.15u W=0.36u AS=0.0684p AD=0.0684p
+ PS=0.74u PD=0.74u
M$25 \$31 \$41 \$42 \$2 sg13_lv_nmos L=0.15u W=0.36u AS=0.0684p AD=0.1224p
+ PS=0.74u PD=1.4u
M$26 \$19 \$8 \$20 \$2 sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.0684p
+ PS=1.4u PD=0.74u
M$27 \$20 \$8 \$23 \$2 sg13_lv_nmos L=0.15u W=0.36u AS=0.0684p AD=0.0684p
+ PS=0.74u PD=0.74u
M$28 \$23 \$8 \$21 \$2 sg13_lv_nmos L=0.15u W=0.36u AS=0.0684p AD=0.0684p
+ PS=0.74u PD=0.74u
M$29 \$21 \$8 \$28 \$2 sg13_lv_nmos L=0.15u W=0.36u AS=0.0684p AD=0.0684p
+ PS=0.74u PD=0.74u
M$30 \$28 \$8 \$17 \$2 sg13_lv_nmos L=0.15u W=0.36u AS=0.0684p AD=0.1224p
+ PS=0.74u PD=1.4u
M$31 \$1 \$41 \$47 \$1 sg13_lv_pmos L=0.15u W=0.32u AS=0.1088p AD=0.0608p
+ PS=1.32u PD=0.7u
M$32 \$47 \$41 \$42 \$1 sg13_lv_pmos L=0.15u W=0.32u AS=0.0608p AD=0.1088p
+ PS=0.7u PD=1.32u
M$33 \$1 \$8 \$4 \$1 sg13_lv_pmos L=0.15u W=0.32u AS=0.1088p AD=0.0608p
+ PS=1.32u PD=0.7u
M$34 \$4 \$8 \$17 \$1 sg13_lv_pmos L=0.15u W=0.32u AS=0.0608p AD=0.1088p
+ PS=0.7u PD=1.32u
M$35 \$8 \$8 \$15 \$1 sg13_lv_pmos L=0.15u W=0.32u AS=0.1088p AD=0.0608p
+ PS=1.32u PD=0.7u
M$36 \$15 \$8 \$7 \$1 sg13_lv_pmos L=0.15u W=0.32u AS=0.0608p AD=0.1088p
+ PS=0.7u PD=1.32u
M$37 \$41 \$41 \$51 \$1 sg13_lv_pmos L=0.15u W=0.32u AS=0.1088p AD=0.0608p
+ PS=1.32u PD=0.7u
M$38 \$51 \$41 \$43 \$1 sg13_lv_pmos L=0.15u W=0.32u AS=0.0608p AD=0.1088p
+ PS=0.7u PD=1.32u
.ENDS PFD
