* Extracted by KLayout with SG13G2 LVS runset on : 01/07/2025 12:53

.SUBCKT charge_pump
M$1 6 5 9 6 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u PD=0.74u
M$2 9 2 8 6 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u PD=1.34u
M$3 6 1 3 6 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u PD=1.34u
M$4 3 1 7 7 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u PD=1.28u
M$5 8 3 10 7 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$6 10 4 7 7 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u PD=1.28u
.ENDS charge_pump
