** sch_path: /foss/designs/Team2/inverter/inverter_tb.sch
**.subckt inverter_tb Vout
*.opin Vout
x1 Vdd Vin Vout GND inverter
Vin Vin GND PULSE(0 1 0.5n 100p 100p 1n 2n)
Vdd Vdd GND 1
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt



.param temp=27
.control
save all
tran 50p 20n
meas tran tdelay TRIG v(Vin) VAL=0.9 FALl=1 TRAG v(Vout) VAl=0.9 RISE=1
write tran_logic_not.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/Team2/inverter/inverter.sym # of pins=4
** sym_path: /foss/designs/Team2/inverter/inverter.sym
** sch_path: /foss/designs/Team2/inverter/inverter.sch
.subckt inverter VP A Y VN
*.iopin VN
*.iopin VP
*.ipin A
*.opin Y
XM1 Y A VP VP sg13_lv_pmos w=2u l=0.13u ng=1 m=1 rfmode=1
XM2 Y A VN VN sg13_lv_nmos w=1u l=0.13u ng=1 m=1 rfmode=1
.ends

.GLOBAL GND
.end
