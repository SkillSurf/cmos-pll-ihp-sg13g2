** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_vco_tb.sch
**.subckt t2_vco_tb Vout
*.opin Vout
VDD net4 GND 1.2
vctl net3 GND 0.8
Ven net2 GND 1.2
Venb net1 GND 0
VNB net5 GND 0
VPB net6 GND 1.2
x1 net4 net6 GND net5 Vout net3 net2 net1 t2_vco
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt



.param temp=27
.ic v(Vout)=0
.tran 10 5u
.save all
.plot v(Vout)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_vco.sym # of pins=8
** sym_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_vco.sym
** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_vco.sch
.subckt t2_vco VPWR VPB VGND VNB Vout vctl en enb
*.iopin VPWR
*.iopin VPB
*.iopin VGND
*.iopin VNB
*.ipin vctl
*.ipin en
*.ipin enb
*.opin Vout
XM1 net1 en VPWR VPB sg13_lv_pmos w=1.0u l=0.15u ng=1 m=1
XM2 net1 net1 VPWR VPB sg13_lv_pmos w=3.0u l=0.15u ng=1 m=1
XM3 vco_source net1 VPWR VPB sg13_lv_pmos w=3.0u l=0.15u ng=1 m=1
XM4 net1 vctl net2 VNB sg13_lv_nmos w=0.75u l=0.15u ng=1 m=2
XM5 net2 net2 VGND VNB sg13_lv_nmos w=1.5u l=0.15u ng=1 m=1
XM6 vco_sink net2 VGND VNB sg13_lv_nmos w=1.5u l=0.15u ng=1 m=1
XM7 net2 enb VGND VNB sg13_lv_nmos w=0.5u l=0.15u ng=1 m=1
XM8 vctl enb VGND VNB sg13_lv_nmos w=0.5u l=0.15u ng=1 m=1
XM9 Vout enb VGND VNB sg13_lv_nmos w=0.5u l=0.15u ng=1 m=1
x1 vco_source VPB Vout net3 VNB vco_sink t2_vco_inverter
x2 vco_source VPB net3 net4 VNB vco_sink t2_vco_inverter
x3 vco_source VPB net4 Vout VNB vco_sink t2_vco_inverter
.ends


* expanding   symbol:  /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_vco_inverter.sym # of pins=6
** sym_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_vco_inverter.sym
** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_vco_inverter.sch
.subckt t2_vco_inverter VPWR VPB A Y VNB VGND
*.iopin VPWR
*.iopin VGND
*.ipin A
*.opin Y
*.iopin VPB
*.iopin VNB
XM2 Y A VPWR VPB sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
XM1 Y A VGND VNB sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
