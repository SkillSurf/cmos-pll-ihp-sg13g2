** sch_path: /foss/designs/Team1/inverter/inverter_tb.sch
**.subckt inverter_tb Vout
*.opin Vout
Vin Vin GND dc 0 ac 0 pulse(0, 1.2, 0, 0.8n, 0.8n, 2n, 4n)
C1 Vout GND 100f m=1
x1 Vout Vin inverter
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt



.param temp=27
.control
save all
tran 50p 20n
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/Team1/inverter/inverter.sym # of pins=2
** sym_path: /foss/designs/Team1/inverter/inverter.sym
** sch_path: /foss/designs/Team1/inverter/inverter.sch
.subckt inverter Y A
*.ipin A
*.opin Y
XM1 Y A net1 net1 sg13_lv_pmos w=2u l=0.13u ng=1 m=1 rfmode=1
XM2 Y A GND GND sg13_lv_nmos w=1u l=0.13u ng=1 m=1 rfmode=1
V1 net1 GND 1.2
.ends

.GLOBAL GND
.end
