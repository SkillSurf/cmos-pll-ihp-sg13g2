* Extracted by KLayout with SG13G2 LVS runset on : 19/07/2025 19:54

.SUBCKT pll_3bitDiv
X$14 \$1 3bit_freq_divider
X$15 \$1 3bit_freq_divider
X$16 \$1 PFD
X$17 \$1 11Stage_vco_new
X$18 \$1 Bias_gen
X$19 \$1 loop_filter
X$20 \$1 charge_pump
X$21 \$I1 \$1 \$I3 \$I4 sg13g2_inv_1
.ENDS pll_3bitDiv

.SUBCKT charge_pump \$9
M$1 \$9 \$5 \$8 \$9 sg13_lv_nmos L=0.13u W=1.2u AS=0.408p AD=0.207p PS=3.08u
+ PD=1.545u
M$2 \$8 \$2 \$7 \$9 sg13_lv_nmos L=0.13u W=1.2u AS=0.207p AD=0.408p PS=1.545u
+ PD=3.08u
M$3 \$7 \$3 \$11 \$6 sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p
+ PS=1.34u PD=0.74u
M$4 \$11 \$4 \$6 \$6 sg13_lv_pmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p
+ PS=0.74u PD=1.34u
M$5 \$3 \$1 \$6 \$6 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
M$6 \$9 \$1 \$3 \$9 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
.ENDS charge_pump

.SUBCKT loop_filter \$1
M$1 \$1 \$4 \$1 \$1 sg13_lv_nmos L=0.65u W=45u AS=9p AD=9p PS=60u PD=60u
R$31 \$4 \$2 rhigh w=0.6u l=0.96u ps=0 b=0 m=1
R$32 \$3 \$4 rhigh w=0.5u l=0.96u ps=0 b=0 m=1
M$33 \$1 \$2 \$1 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.201p AD=0.201p PS=2.68u
+ PD=2.68u
M$35 \$1 \$3 \$1 \$1 sg13_lv_nmos L=0.65u W=15u AS=3p AD=3p PS=28u PD=28u
.ENDS loop_filter

.SUBCKT Bias_gen \$1
R$1 \$11 \$13 rhigh w=1u l=12u ps=0 b=0 m=1
R$2 \$3 \$2 rhigh w=1u l=12u ps=0 b=0 m=1
M$3 \$10 \$6 \$2 \$1 sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$4 \$8 \$6 \$3 \$1 sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$5 \$6 \$6 \$2 \$1 sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$6 \$8 \$10 \$7 \$1 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$7 \$6 \$4 \$2 \$1 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$8 \$7 \$5 \$2 \$1 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$9 \$6 \$8 \$11 \$9 sg13_lv_pmos L=1u W=4u AS=1.06p AD=1.06p PS=7.06u PD=7.06u
M$11 \$13 \$8 \$8 \$9 sg13_lv_pmos L=1u W=2u AS=0.68p AD=0.68p PS=4.68u PD=4.68u
M$12 \$13 \$12 \$12 \$9 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$13 \$13 \$5 \$8 \$9 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$14 \$12 \$10 \$10 \$9 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$15 \$13 \$5 \$10 \$9 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
.ENDS Bias_gen

.SUBCKT 11Stage_vco_new VGND
M$1 \$83 \$61 \$52 VGND sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u
+ PD=2.62u
M$3 VGND vctl \$137 VGND sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p
+ PS=2.02u PD=2.02u
M$5 VGND vctl \$142 VGND sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p
+ PS=2.02u PD=2.02u
M$7 \$86 \$35 \$71 VGND sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u
+ PD=2.62u
M$9 \$84 \$68 \$61 VGND sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u
+ PD=2.62u
M$11 VGND vctl \$84 VGND sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p
+ PS=2.02u PD=2.02u
M$13 VGND vctl \$126 VGND sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p
+ PS=2.02u PD=2.02u
M$15 \$87 \$81 \$35 VGND sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u
+ PD=2.62u
M$17 VGND vctl \$36 VGND sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p
+ PS=2.02u PD=2.02u
M$19 \$85 \$71 \$68 VGND sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u
+ PD=2.62u
M$21 VGND vctl \$85 VGND sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p
+ PS=2.02u PD=2.02u
M$23 VGND vctl \$125 VGND sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p
+ PS=2.02u PD=2.02u
M$25 VGND vctl \$132 VGND sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p
+ PS=2.02u PD=2.02u
M$27 VGND vctl \$87 VGND sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p
+ PS=2.02u PD=2.02u
M$29 VGND vctl \$82 VGND sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p
+ PS=2.02u PD=2.02u
M$31 VGND vctl \$86 VGND sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p
+ PS=2.02u PD=2.02u
M$33 \$82 \$52 \$46 VGND sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u
+ PD=2.62u
M$35 VGND vctl \$83 VGND sg13_lv_nmos L=0.13u W=0.6u AS=0.168p AD=0.168p
+ PS=2.02u PD=2.02u
M$37 \$25 \$36 VPWR VPWR sg13_lv_pmos L=0.13u W=0.8u AS=0.2825p AD=0.281p
+ PS=3.57u PD=3.56u
M$41 \$152 \$36 VPWR VPWR sg13_lv_pmos L=0.13u W=0.8u AS=0.2375p AD=0.326p
+ PS=2.97u PD=4.16u
M$45 \$153 \$36 VPWR VPWR sg13_lv_pmos L=0.13u W=0.8u AS=0.2375p AD=0.326p
+ PS=2.97u PD=4.16u
M$49 \$3 \$36 VPWR VPWR sg13_lv_pmos L=0.13u W=0.8u AS=0.2825p AD=0.281p
+ PS=3.57u PD=3.56u
M$53 \$4 \$36 VPWR VPWR sg13_lv_pmos L=0.13u W=0.8u AS=0.2825p AD=0.281p
+ PS=3.57u PD=3.56u
M$57 \$35 \$81 \$7 VPWR sg13_lv_pmos L=0.13u W=2u AS=0.5012p AD=0.5p PS=4.51u
+ PD=4.5u
M$61 \$46 \$52 \$3 VPWR sg13_lv_pmos L=0.13u W=2u AS=0.5012p AD=0.5p PS=4.51u
+ PD=4.5u
M$65 \$31 \$36 VPWR VPWR sg13_lv_pmos L=0.13u W=0.8u AS=0.2825p AD=0.281p
+ PS=3.57u PD=3.56u
M$69 \$68 \$71 \$31 VPWR sg13_lv_pmos L=0.13u W=2u AS=0.5012p AD=0.5p PS=4.51u
+ PD=4.5u
M$73 \$7 \$36 VPWR VPWR sg13_lv_pmos L=0.13u W=0.8u AS=0.2825p AD=0.281p
+ PS=3.57u PD=3.56u
M$77 VPWR \$36 \$36 VPWR sg13_lv_pmos L=0.13u W=0.8u AS=0.28175p AD=0.28175p
+ PS=3.565u PD=3.565u
M$81 \$18 \$36 VPWR VPWR sg13_lv_pmos L=0.13u W=0.8u AS=0.2825p AD=0.281p
+ PS=3.57u PD=3.56u
M$85 \$61 \$68 \$25 VPWR sg13_lv_pmos L=0.13u W=2u AS=0.5012p AD=0.5p PS=4.51u
+ PD=4.5u
M$89 \$155 \$36 VPWR VPWR sg13_lv_pmos L=0.13u W=0.8u AS=0.2375p AD=0.326p
+ PS=2.97u PD=4.16u
M$93 \$71 \$35 \$18 VPWR sg13_lv_pmos L=0.13u W=2u AS=0.5012p AD=0.5p PS=4.51u
+ PD=4.5u
M$97 \$151 \$36 VPWR VPWR sg13_lv_pmos L=0.13u W=0.8u AS=0.2375p AD=0.326p
+ PS=2.97u PD=4.16u
M$101 \$52 \$61 \$4 VPWR sg13_lv_pmos L=0.13u W=2u AS=0.5012p AD=0.5p PS=4.51u
+ PD=4.5u
M$105 \$154 \$36 VPWR VPWR sg13_lv_pmos L=0.13u W=0.8u AS=0.2375p AD=0.326p
+ PS=2.97u PD=4.16u
M$109 VGND \$81 Vout VGND sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u
+ PD=2.62u
M$111 VPWR \$81 Vout VPWR sg13_lv_pmos L=0.13u W=2u AS=0.5p AD=0.5p PS=4.5u
+ PD=4.5u
C$115 VGND \$81 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$116 VGND \$35 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$117 VGND \$129 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$118 VGND \$127 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$119 VGND \$46 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$120 VGND \$148 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$121 VGND \$71 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$122 VGND \$128 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$123 VGND Vout cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=2
C$124 VGND \$61 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$125 VGND \$68 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$127 VGND \$52 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
M$128 \$132 \$46 \$127 VGND sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p
+ PS=2.62u PD=2.62u
M$130 \$127 \$46 \$151 VPWR sg13_lv_pmos L=0.13u W=2u AS=0.4412p AD=0.56p
+ PS=3.77u PD=5.24u
M$134 \$137 \$127 \$128 VGND sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p
+ PS=2.62u PD=2.62u
M$136 \$128 \$127 \$152 VPWR sg13_lv_pmos L=0.13u W=2u AS=0.4412p AD=0.56p
+ PS=3.77u PD=5.24u
M$140 \$142 \$128 \$148 VGND sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p
+ PS=2.62u PD=2.62u
M$142 \$148 \$128 \$153 VPWR sg13_lv_pmos L=0.13u W=2u AS=0.4412p AD=0.56p
+ PS=3.77u PD=5.24u
M$146 \$125 \$148 \$129 VGND sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p
+ PS=2.62u PD=2.62u
M$148 \$129 \$148 \$154 VPWR sg13_lv_pmos L=0.13u W=2u AS=0.4412p AD=0.56p
+ PS=3.77u PD=5.24u
M$152 \$126 \$129 \$81 VGND sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p
+ PS=2.62u PD=2.62u
M$154 \$81 \$129 \$155 VPWR sg13_lv_pmos L=0.13u W=2u AS=0.4412p AD=0.56p
+ PS=3.77u PD=5.24u
.ENDS 11Stage_vco_new

.SUBCKT PFD VSS
M$1 \$5 VCO_CLK \$7 VSS sg13_lv_nmos L=0.15u W=0.84u AS=0.2226p AD=0.2226p
+ PS=2.32u PD=2.32u
M$3 \$10 Ref_CLK \$12 VSS sg13_lv_nmos L=0.15u W=0.84u AS=0.2226p AD=0.2226p
+ PS=2.32u PD=2.32u
M$5 VSS \$13 UP VSS sg13_lv_nmos L=0.15u W=0.48u AS=0.1632p AD=0.1632p PS=1.64u
+ PD=1.64u
M$6 VSS \$4 DOWN VSS sg13_lv_nmos L=0.15u W=0.48u AS=0.1632p AD=0.1632p
+ PS=1.64u PD=1.64u
M$7 \$9 VCO_CLK VSS VSS sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p
+ PS=1.4u PD=1.4u
M$8 VSS \$10 \$13 VSS sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p
+ PS=1.4u PD=1.4u
M$9 VSS \$5 \$4 VSS sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p PS=1.4u
+ PD=1.4u
M$10 \$8 Ref_CLK VSS VSS sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p
+ PS=1.4u PD=1.4u
M$11 VDD \$13 UP VDD sg13_lv_pmos L=0.15u W=0.96u AS=0.2304p AD=0.2304p
+ PS=2.72u PD=2.72u
M$14 VDD \$4 DOWN VDD sg13_lv_pmos L=0.15u W=0.96u AS=0.2304p AD=0.2304p
+ PS=2.72u PD=2.72u
M$17 \$13 \$10 VDD VDD sg13_lv_pmos L=0.15u W=0.72u AS=0.1908p AD=0.1908p
+ PS=2.14u PD=2.14u
M$19 VDD \$5 \$4 VDD sg13_lv_pmos L=0.15u W=0.72u AS=0.1908p AD=0.1908p
+ PS=2.14u PD=2.14u
M$21 \$9 Ref_CLK \$12 VSS sg13_lv_nmos L=0.15u W=1.8u AS=0.396p AD=0.396p
+ PS=4.36u PD=4.36u
M$26 \$8 VCO_CLK \$7 VSS sg13_lv_nmos L=0.15u W=1.8u AS=0.396p AD=0.396p
+ PS=4.36u PD=4.36u
M$31 \$12 Ref_CLK VDD VDD sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p AD=0.1696p
+ PS=2.02u PD=2.02u
M$33 \$7 VCO_CLK VDD VDD sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p AD=0.1696p
+ PS=2.02u PD=2.02u
M$35 \$5 VCO_CLK VCO_CLK VDD sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p AD=0.1696p
+ PS=2.02u PD=2.02u
M$37 \$10 Ref_CLK Ref_CLK VDD sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p
+ AD=0.1696p PS=2.02u PD=2.02u
.ENDS PFD

.SUBCKT 3bit_freq_divider VSS
X$1 \$17 VDD VSS sg13g2_tiehi
X$2 \$8 \$13 \$13 CLK_OUT VSS \$17 VDD dff_nclk
X$3 VDD VSS \$10 \$11 \$9 \$8 sg13g2_or3_1
X$4 \$22 \$18 \$5 A1 \$9 VSS \$8 VDD freq_div_cell
X$5 \$29 \$22 \$5 A0 \$10 VSS \$8 VDD freq_div_cell
X$6 \$29 VDD VSS sg13g2_tiehi
X$7 \$18 \$I25 \$5 A2 \$11 VSS \$8 VDD freq_div_cell
X$8 VDD VSS \$5 CLK_IN EN sg13g2_nand2_1
.ENDS 3bit_freq_divider

.SUBCKT sg13g2_nand2_1 VDD VSS Y A B
M$1 VSS B \$6 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.0666p PS=2.16u
+ PD=0.92u
M$2 \$6 A Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.0666p AD=0.2516p PS=0.92u
+ PD=2.16u
M$3 VDD B Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.2128p PS=2.92u
+ PD=1.5u
M$4 Y A VDD VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.3808p PS=1.5u
+ PD=2.92u
.ENDS sg13g2_nand2_1

.SUBCKT sg13g2_or3_1 VDD VSS C A B X
M$1 \$6 C VSS VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.187p AD=0.1045p PS=1.78u
+ PD=0.93u
M$2 VSS B \$6 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.1045p AD=0.198p PS=0.93u
+ PD=1.27u
M$3 \$6 A VSS VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.198p AD=0.13395p PS=1.27u
+ PD=1.12u
M$4 VSS \$6 X VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.13395p AD=0.2516p PS=1.12u
+ PD=2.16u
M$5 \$6 C \$9 VDD sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.1275p PS=2.68u
+ PD=1.255u
M$6 \$9 B \$8 VDD sg13_lv_pmos L=0.13u W=1u AS=0.1275p AD=0.22p PS=1.255u
+ PD=1.44u
M$7 \$8 A VDD VDD sg13_lv_pmos L=0.13u W=1u AS=0.22p AD=0.3822p PS=1.44u
+ PD=1.84u
M$8 VDD \$6 X VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3822p AD=0.3808p PS=1.84u
+ PD=2.92u
.ENDS sg13g2_or3_1

.SUBCKT sg13g2_tiehi L_HI VDD VSS
M$1 VSS \$4 \$4 VSS sg13_lv_nmos L=0.13u W=0.3u AS=0.2307p AD=0.102p PS=1.615u
+ PD=1.28u
M$2 VSS \$3 \$1 VSS sg13_lv_nmos L=0.13u W=0.795u AS=0.2307p AD=0.274275p
+ PS=1.615u PD=2.28u
M$3 \$3 \$4 VDD VDD sg13_lv_pmos L=0.13u W=0.66u AS=0.2442p AD=0.4657125p
+ PS=2.06u PD=2.54u
M$4 VDD \$1 L_HI VDD sg13_lv_pmos L=0.13u W=1.155u AS=0.4657125p AD=0.3927p
+ PS=2.54u PD=2.99u
.ENDS sg13g2_tiehi

.SUBCKT freq_div_cell Cin Cout CLK BIT DIV \$7 nRST \$11
X$1 Cin \$6 \$9 Cout \$7 \$11 half_add
X$2 CLK \$9 \$I8 \$6 \$7 nRST \$11 dff_nclk
X$3 \$7 DIV \$11 \$6 BIT sg13g2_xor2_1
.ENDS freq_div_cell

.SUBCKT dff_nclk nCLK D nQ Q \$6 nRST \$9
X$1 \$9 \$6 nCLK \$5 sg13g2_inv_1
X$2 \$6 nRST nQ Q D \$5 \$9 sg13g2_dfrbp_1
.ENDS dff_nclk

.SUBCKT half_add inA inB sum cout \$5 \$6
X$1 \$5 sum \$6 inA inB sg13g2_xor2_1
X$2 \$6 \$5 cout inA inB sg13g2_and2_1
.ENDS half_add

.SUBCKT sg13g2_dfrbp_1 VSS RESET_B Q_N Q D CLK VDD
M$1 \$8 \$5 VSS VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.187p AD=0.14505p PS=1.78u
+ PD=1.15u
M$2 VSS \$8 Q VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.14505p AD=0.2516p PS=1.15u
+ PD=2.16u
M$3 \$4 D \$15 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.0504p PS=1.52u
+ PD=0.66u
M$4 \$15 RESET_B VSS VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.0504p AD=0.1428p
+ PS=0.66u PD=1.52u
M$5 \$5 \$11 \$19 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.2017p AD=0.0546p
+ PS=1.48u PD=0.68u
M$6 \$19 \$6 VSS VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.0546p AD=0.0903p
+ PS=0.68u PD=0.85u
M$7 VSS RESET_B \$18 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.0903p AD=0.04725p
+ PS=0.85u PD=0.645u
M$8 \$18 \$5 \$6 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.04725p AD=0.1428p
+ PS=0.645u PD=1.52u
M$9 VSS \$13 \$14 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.1825p AD=0.193975p
+ PS=1.325u PD=1.29u
M$10 \$14 \$3 \$5 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.193975p AD=0.2017p
+ PS=1.29u PD=1.48u
M$11 \$4 \$11 \$13 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p
+ PS=1.52u PD=0.8u
M$12 \$13 \$3 \$16 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.0798p AD=0.0546p
+ PS=0.8u PD=0.68u
M$13 \$16 \$14 \$17 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.0546p AD=0.0483p
+ PS=0.68u PD=0.65u
M$14 VSS RESET_B \$17 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1825p AD=0.0483p
+ PS=1.325u PD=0.65u
M$15 VSS CLK \$11 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1544p AD=0.2516p
+ PS=1.235u PD=2.16u
M$16 VSS \$11 \$3 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1544p AD=0.2516p
+ PS=1.235u PD=2.16u
M$17 VSS \$5 Q_N VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.2775p
+ PS=2.16u PD=2.23u
M$18 \$11 CLK VDD VDD sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.19p PS=2.68u
+ PD=1.38u
M$19 VDD \$11 \$3 VDD sg13_lv_pmos L=0.13u W=1u AS=0.19p AD=0.34p PS=1.38u
+ PD=2.68u
M$20 VDD D \$4 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p PS=1.52u
+ PD=0.8u
M$21 \$4 RESET_B VDD VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.1428p
+ PS=0.8u PD=1.52u
M$22 VDD \$5 \$8 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2016p AD=0.2856p PS=1.5u
+ PD=2.36u
M$23 VDD \$8 Q VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2016p AD=0.3808p PS=1.5u
+ PD=2.92u
M$24 VDD \$13 \$14 VDD sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.19p PS=2.68u
+ PD=1.38u
M$25 \$14 \$11 \$5 VDD sg13_lv_pmos L=0.13u W=1u AS=0.19p AD=0.17695p PS=1.38u
+ PD=1.56u
M$26 \$5 \$3 \$22 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.17695p AD=0.04305p
+ PS=1.56u PD=0.625u
M$27 \$22 \$6 VDD VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.04305p AD=0.0798p
+ PS=0.625u PD=0.8u
M$28 VDD RESET_B \$6 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.0798p
+ PS=0.8u PD=0.8u
M$29 VDD \$5 \$6 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.2163p AD=0.0798p
+ PS=1.55u PD=0.8u
M$30 VDD \$5 Q_N VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2163p AD=0.7616p
+ PS=1.55u PD=3.6u
M$31 \$4 \$3 \$13 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p
+ PS=1.52u PD=0.8u
M$32 \$13 \$11 \$21 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.05145p
+ PS=0.8u PD=0.665u
M$33 \$21 \$14 VDD VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.05145p AD=0.11785p
+ PS=0.665u PD=1.025u
M$34 VDD RESET_B \$13 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.11785p AD=0.1533p
+ PS=1.025u PD=1.57u
.ENDS sg13g2_dfrbp_1

.SUBCKT sg13g2_inv_1 VDD VSS A Y
M$1 VSS A Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p AD=0.259p PS=2.18u
+ PD=2.18u
M$2 VDD A Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p AD=0.392p PS=2.94u
+ PD=2.94u
.ENDS sg13g2_inv_1

.SUBCKT sg13g2_and2_1 VDD VSS X A B
M$1 \$6 A \$7 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.2176p AD=0.1216p PS=1.96u
+ PD=1.02u
M$2 VSS B \$7 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.1331p AD=0.1216p PS=1.12u
+ PD=1.02u
M$3 VSS \$6 X VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1331p AD=0.2516p PS=1.12u
+ PD=2.16u
M$4 VDD A \$6 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p AD=0.1596p PS=2.36u
+ PD=1.22u
M$5 VDD B \$6 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.1918p AD=0.1596p PS=1.5u
+ PD=1.22u
M$6 VDD \$6 X VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.1918p AD=0.3808p PS=1.5u
+ PD=2.92u
.ENDS sg13g2_and2_1

.SUBCKT sg13g2_xor2_1 VSS X VDD A B
M$1 VSS A \$1 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.374p AD=0.174625p PS=2.46u
+ PD=1.185u
M$2 VSS B \$1 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.15245p AD=0.174625p
+ PS=1.17u PD=1.185u
M$3 VSS A \$8 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.15245p AD=0.0888p PS=1.17u
+ PD=0.98u
M$4 \$8 B X VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.0888p AD=0.1628p PS=0.98u
+ PD=1.18u
M$5 X \$1 VSS VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1628p AD=0.3108p PS=1.18u
+ PD=2.32u
M$6 \$3 A VDD VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.2128p PS=2.92u
+ PD=1.5u
M$7 VDD B \$3 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.2128p PS=1.5u
+ PD=1.5u
M$8 \$3 \$1 X VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.3808p PS=1.5u
+ PD=2.92u
M$9 VDD A \$9 VDD sg13_lv_pmos L=0.13u W=1u AS=0.36p AD=0.1225p PS=2.72u
+ PD=1.245u
M$10 \$9 B \$1 VDD sg13_lv_pmos L=0.13u W=1u AS=0.1225p AD=0.34p PS=1.245u
+ PD=2.68u
.ENDS sg13g2_xor2_1
