** sch_path: /foss/designs/iic-osic-tools/cmos-pll-ihp-sg13g2/Combined_Design/design_data/xschem/pll_3bitDiv_tb.sch

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ_stat
.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ
.include /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice

**.subckt pll_3bitDiv_tb
V1 VDD GND 1.2
V2 CLK_IN GND PULSE(0 1.2 0.2n 5n 5n 50n 100n)
Va0 A0 GND dc {A0}
Va1 A1 GND dc {A1}
* noconn CLK_OUT
Va2 A2 GND dc {A2}
Vb0 B0 GND dc {B0}
Vb1 B1 GND dc {B1}
Vb2 B2 GND dc {B2}
x1 CLK_IN CLK_OUT B0 B2 B1 VDD GND GND A1 A2 A0 pll_3bitDiv
**** begin user architecture code


.include pll_3bitDiv.pex.spice
.param temp=27
.options method=gear
.options gmin=1e-10

.control
save all

tran 1n 1u uic

write tran_pll_3bitDiv_tb_post.raw
.endc





.param A0 = 1.2
.param A1 = 0
.param A2 = 0




.param B0 = 1.2
.param B1 = 0
.param B2 = 0


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
