* NGSPICE file created from 11Stage_vco_new_update2.ext - technology: ihp-sg13g2

.subckt x11Stage_vco_new_update2 vctl VPWR VGND Vout
X0 a_542_269# a_745_n2395# a_684_n1958# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X1 a_7398_n1956# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X2 a_4776_351# a_3434_351# a_4909_n217# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X3 a_4909_n217# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X4 Vout a_7212_321# VPWR VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X5 a_4771_n2395# a_6113_n2395# a_6051_n2525# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X6 a_2026_n1958# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X7 a_6024_351# a_4776_351# a_6118_351# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X8 a_4909_n217# a_3434_351# a_4776_351# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X9 a_6113_n2395# a_6118_351# a_7397_n2523# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X10 a_656_351# a_542_269# a_750_351# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X11 a_7397_n2523# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X12 VGND vctl a_4909_n217# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X13 a_3434_351# VGND cap_cmim l=6.99u w=6.99u
X14 VPWR a_7212_321# Vout VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X15 VPWR a_620_930# a_3367_n2525# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X16 a_3340_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X17 a_2092_351# a_750_351# a_1998_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X18 a_6051_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X19 VPWR a_620_930# a_3367_n2525# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X20 a_684_n1958# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X21 VPWR a_620_930# a_4682_351# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X22 a_683_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X23 a_6052_n1958# a_6113_n2395# a_4771_n2395# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X24 a_2092_351# a_750_351# a_1998_351# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X25 a_7398_n1956# a_6118_351# a_6113_n2395# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X26 VPWR a_620_930# a_3340_351# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X27 VGND a_7198_n376# Vout VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X28 a_7397_n2523# a_6118_351# a_6113_n2395# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X29 a_2025_n2525# a_2087_n2395# a_745_n2395# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X30 VPWR a_620_930# a_4709_n2525# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X31 a_4709_n2525# a_4771_n2395# a_3429_n2395# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X32 VPWR a_620_930# a_2025_n2525# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X33 a_2025_n2525# a_2087_n2395# a_745_n2395# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X34 VGND vctl a_6052_n1958# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X35 VGND vctl a_7398_n1956# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X36 Vout a_7212_321# VPWR VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X37 a_6251_n217# a_4776_351# a_6118_351# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X38 VPWR a_620_930# a_7397_n2523# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X39 VGND vctl a_6251_n217# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X40 VPWR a_7212_321# Vout VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X41 a_883_n217# a_542_269# a_750_351# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X42 VGND vctl a_883_n217# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X43 VPWR a_620_930# a_3340_351# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X44 a_2092_351# a_750_351# a_2225_n217# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X45 a_2225_n217# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X46 a_3367_n2525# a_3429_n2395# a_2087_n2395# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X47 a_4682_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X48 Vout VGND cap_cmim l=6.99u w=6.99u
X49 a_4771_n2395# a_6113_n2395# a_6051_n2525# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X50 a_3367_n2525# a_3429_n2395# a_2087_n2395# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X51 a_6024_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X52 a_6113_n2395# a_6118_351# a_7397_n2523# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X53 a_542_269# a_745_n2395# a_683_n2525# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X54 a_3340_351# a_2092_351# a_3434_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X55 a_2025_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X56 a_745_n2395# a_2087_n2395# a_2025_n2525# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X57 a_1998_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X58 a_542_269# VGND cap_cmim l=6.99u w=6.99u
X59 a_2025_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X60 a_656_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X61 a_745_n2395# a_2087_n2395# a_2025_n2525# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X62 a_683_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X63 a_620_930# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X64 a_2087_n2395# a_3429_n2395# a_3368_n1958# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X65 a_542_269# a_745_n2395# a_683_n2525# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X66 VPWR a_620_930# a_4709_n2525# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X67 VPWR a_620_930# a_6024_351# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X68 a_684_n1958# a_745_n2395# a_542_269# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X69 a_1998_351# a_750_351# a_2092_351# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X70 VPWR a_620_930# a_656_351# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X71 a_2225_n217# a_750_351# a_2092_351# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X72 VGND vctl a_2225_n217# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X73 VPWR a_620_930# a_620_930# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X74 a_3368_n1958# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X75 a_3429_n2395# VGND cap_cmim l=6.99u w=6.99u
X76 a_3434_351# a_2092_351# a_3340_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X77 a_3367_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X78 a_4682_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X79 a_3434_351# a_2092_351# a_3567_n217# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X80 a_3567_n217# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X81 a_620_930# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X82 a_2087_n2395# a_3429_n2395# a_3367_n2525# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X83 VPWR a_620_930# a_6051_n2525# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X84 a_3429_n2395# a_4771_n2395# a_4710_n1958# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X85 VGND vctl a_684_n1958# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X86 a_4682_351# a_3434_351# a_4776_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X87 a_4771_n2395# VGND cap_cmim l=6.99u w=6.99u
X88 a_6051_n2525# a_6113_n2395# a_4771_n2395# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X89 a_6118_351# a_4776_351# a_6251_n217# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X90 a_6251_n217# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X91 VPWR a_620_930# a_6024_351# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X92 VPWR a_620_930# a_6051_n2525# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X93 a_6051_n2525# a_6113_n2395# a_4771_n2395# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X94 a_3434_351# a_2092_351# a_3340_351# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X95 a_4682_351# a_3434_351# a_4776_351# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X96 VPWR a_620_930# a_656_351# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X97 a_6118_351# VGND cap_cmim l=6.99u w=6.99u
X98 a_4710_n1958# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X99 a_3368_n1958# a_3429_n2395# a_2087_n2395# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X100 a_3340_351# a_2092_351# a_3434_351# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X101 a_4709_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X102 a_4771_n2395# a_6113_n2395# a_6052_n1958# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X103 a_656_351# a_542_269# a_750_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X104 a_2087_n2395# VGND cap_cmim l=6.99u w=6.99u
X105 VGND vctl a_620_930# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X106 a_6118_351# a_4776_351# a_6024_351# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X107 a_2092_351# VGND cap_cmim l=6.99u w=6.99u
X108 a_4709_n2525# a_4771_n2395# a_3429_n2395# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X109 VPWR a_620_930# a_620_930# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X110 a_4776_351# a_3434_351# a_4682_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X111 a_750_351# VGND cap_cmim l=6.99u w=6.99u
X112 VGND vctl a_3368_n1958# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X113 a_4709_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X114 VPWR a_620_930# a_683_n2525# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X115 a_7397_n2523# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X116 a_683_n2525# a_745_n2395# a_542_269# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X117 a_4776_351# a_3434_351# a_4682_351# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X118 a_6052_n1958# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X119 a_6113_n2395# VGND cap_cmim l=6.99u w=6.99u
X120 a_620_930# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X121 a_2026_n1958# a_2087_n2395# a_745_n2395# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X122 a_6024_351# a_4776_351# a_6118_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X123 a_6051_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X124 a_4710_n1958# a_4771_n2395# a_3429_n2395# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X125 a_745_n2395# VGND cap_cmim l=6.99u w=6.99u
X126 a_750_351# a_542_269# a_656_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X127 a_4776_351# VGND cap_cmim l=6.99u w=6.99u
X128 VPWR a_620_930# a_1998_351# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X129 a_7397_n2523# a_6118_351# a_6113_n2395# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X130 VGND vctl a_2026_n1958# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X131 a_1998_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X132 a_3367_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X133 a_2087_n2395# a_3429_n2395# a_3367_n2525# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X134 VGND vctl a_4710_n1958# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X135 a_3340_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X136 a_750_351# a_542_269# a_656_351# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X137 a_750_351# a_542_269# a_883_n217# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X138 a_883_n217# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X139 a_6118_351# a_4776_351# a_6024_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X140 VPWR a_620_930# a_4682_351# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X141 a_6024_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X142 VPWR a_620_930# a_683_n2525# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X143 a_3429_n2395# a_4771_n2395# a_4709_n2525# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X144 a_683_n2525# a_745_n2395# a_542_269# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X145 Vout a_7198_n376# VGND VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X146 a_1998_351# a_750_351# a_2092_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X147 a_6113_n2395# a_6118_351# a_7398_n1956# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X148 a_656_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X149 VPWR a_620_930# a_7397_n2523# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X150 VPWR a_620_930# a_2025_n2525# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X151 VPWR a_620_930# a_1998_351# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X152 a_745_n2395# a_2087_n2395# a_2026_n1958# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X153 Vout VGND cap_cmim l=6.99u w=6.99u
X154 a_3567_n217# a_2092_351# a_3434_351# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X155 VGND vctl a_3567_n217# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X156 a_3429_n2395# a_4771_n2395# a_4709_n2525# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
C0 vctl a_3434_351# 0.02497f
C1 a_3340_351# a_3434_351# 0.42148f
C2 a_4682_351# a_3434_351# 0.09926f
C3 a_4776_351# a_4909_n217# 0.22378f
C4 VPWR a_2225_n217# 0.01623f
C5 a_620_930# a_4709_n2525# 0.18962f
C6 a_3429_n2395# a_4710_n1958# 0.23035f
C7 a_6024_351# a_6118_351# 0.4131f
C8 a_745_n2395# a_683_n2525# 0.10818f
C9 a_745_n2395# vctl 0.04038f
C10 a_4776_351# a_620_930# 0.04298f
C11 a_6113_n2395# a_6118_351# 0.81343f
C12 vctl a_6118_351# 0.20887f
C13 a_7198_n376# Vout 0.01195f
C14 a_4771_n2395# a_620_930# 0.04406f
C15 a_7397_n2523# a_6113_n2395# 0.46077f
C16 vctl a_2026_n1958# 0.04894f
C17 a_6052_n1958# a_6118_351# 0.02056f
C18 a_750_351# a_2225_n217# 0.03153f
C19 vctl a_3567_n217# 0.0811f
C20 Vout a_6118_351# 0.77478f
C21 a_745_n2395# a_684_n1958# 0.04971f
C22 VPWR a_6051_n2525# 1.38336f
C23 a_3368_n1958# VPWR 0.01475f
C24 a_2225_n217# a_2092_351# 0.22378f
C25 a_3368_n1958# a_3429_n2395# 0.03778f
C26 a_4771_n2395# a_4709_n2525# 0.11922f
C27 vctl a_6113_n2395# 0.02267f
C28 a_745_n2395# a_2025_n2525# 0.42019f
C29 a_6051_n2525# a_620_930# 0.19288f
C30 a_6052_n1958# a_6113_n2395# 0.03243f
C31 vctl a_6052_n1958# 0.04998f
C32 VPWR a_3434_351# 1.00449f
C33 vctl Vout 0.02121f
C34 a_7398_n1956# a_6118_351# 0.12881f
C35 a_4771_n2395# a_4710_n1958# 0.03159f
C36 vctl a_684_n1958# 0.04284f
C37 a_6251_n217# a_6118_351# 0.2448f
C38 vctl a_883_n217# 0.08086f
C39 a_745_n2395# VPWR 0.81739f
C40 a_3368_n1958# a_2087_n2395# 0.23444f
C41 VPWR a_6118_351# 1.28569f
C42 a_3434_351# a_4909_n217# 0.03153f
C43 a_3367_n2525# VPWR 1.37334f
C44 a_3367_n2525# a_3429_n2395# 0.12854f
C45 a_745_n2395# a_542_269# 0.40206f
C46 a_3434_351# a_620_930# 0.04103f
C47 a_7397_n2523# VPWR 1.38295f
C48 VPWR a_2026_n1958# 0.01457f
C49 a_7212_321# a_6118_351# 0.02041f
C50 VPWR a_3567_n217# 0.0108f
C51 a_7398_n1956# a_6113_n2395# 0.21632f
C52 vctl a_7398_n1956# 0.05123f
C53 a_6051_n2525# a_4771_n2395# 0.46167f
C54 a_745_n2395# a_620_930# 0.08011f
C55 a_620_930# a_6118_351# 0.16863f
C56 a_3434_351# a_2092_351# 0.88103f
C57 vctl a_6251_n217# 0.08336f
C58 a_6024_351# VPWR 1.37111f
C59 a_3367_n2525# a_620_930# 0.19098f
C60 VPWR a_683_n2525# 1.35573f
C61 vctl VPWR 0.28629f
C62 VPWR a_6113_n2395# 1.36426f
C63 a_3429_n2395# vctl 0.04109f
C64 a_3340_351# VPWR 1.36686f
C65 a_4682_351# VPWR 1.35049f
C66 a_7397_n2523# a_620_930# 0.19389f
C67 a_2087_n2395# a_745_n2395# 0.35714f
C68 a_542_269# a_683_n2525# 0.45412f
C69 a_3367_n2525# a_2087_n2395# 0.45379f
C70 a_4776_351# a_3434_351# 0.91818f
C71 vctl a_4909_n217# 0.08436f
C72 a_2087_n2395# a_2026_n1958# 0.03943f
C73 a_6024_351# a_620_930# 0.10045f
C74 VPWR Vout 0.79524f
C75 a_683_n2525# a_620_930# 0.23019f
C76 a_4776_351# a_6118_351# 0.20869f
C77 a_3567_n217# a_2092_351# 0.03153f
C78 a_620_930# a_6113_n2395# 0.06975f
C79 vctl a_620_930# 0.09057f
C80 a_3340_351# a_620_930# 0.19603f
C81 a_4682_351# a_620_930# 0.19696f
C82 a_750_351# vctl 0.02282f
C83 a_542_269# a_684_n1958# 0.23665f
C84 Vout a_7212_321# 0.09147f
C85 a_2087_n2395# a_683_n2525# 0.01232f
C86 a_542_269# a_883_n217# 0.03491f
C87 a_2087_n2395# vctl 0.04184f
C88 vctl a_2092_351# 0.0248f
C89 a_3340_351# a_2092_351# 0.10275f
C90 a_2025_n2525# VPWR 1.36925f
C91 VPWR a_1998_351# 1.37065f
C92 a_684_n1958# a_620_930# 0.06371f
C93 a_6024_351# a_4776_351# 0.1057f
C94 a_883_n217# a_620_930# 0.02036f
C95 vctl a_4776_351# 0.026f
C96 a_4682_351# a_4776_351# 0.42665f
C97 a_750_351# a_883_n217# 0.22378f
C98 a_4771_n2395# a_6113_n2395# 0.58365f
C99 vctl a_4771_n2395# 0.03129f
C100 a_3429_n2395# VPWR 1.08631f
C101 a_2025_n2525# a_620_930# 0.18981f
C102 a_1998_351# a_620_930# 0.19723f
C103 vctl a_2225_n217# 0.07714f
C104 vctl a_4710_n1958# 0.05026f
C105 a_542_269# VPWR 0.7984f
C106 a_750_351# a_1998_351# 0.09188f
C107 Vout a_4776_351# 0.18866f
C108 a_7398_n1956# a_620_930# 0.01439f
C109 a_4771_n2395# a_6052_n1958# 0.22936f
C110 a_2087_n2395# a_2025_n2525# 0.12991f
C111 VPWR a_7212_321# 0.44048f
C112 a_2092_351# a_1998_351# 0.42202f
C113 VPWR a_620_930# 13.1884f
C114 a_3429_n2395# a_620_930# 0.04637f
C115 a_750_351# VPWR 1.05125f
C116 VPWR a_656_351# 1.37421f
C117 a_542_269# a_620_930# 0.93638f
C118 a_7198_n376# a_6118_351# 0.01604f
C119 a_750_351# a_542_269# 0.3548f
C120 a_2087_n2395# VPWR 1.15543f
C121 a_542_269# a_656_351# 0.08875f
C122 a_2087_n2395# a_3429_n2395# 0.72984f
C123 VPWR a_2092_351# 1.29553f
C124 a_6051_n2525# a_6113_n2395# 0.10827f
C125 a_3368_n1958# vctl 0.05041f
C126 VPWR a_4709_n2525# 1.36202f
C127 a_3429_n2395# a_4709_n2525# 0.45955f
C128 a_4776_351# a_6251_n217# 0.03205f
C129 a_750_351# a_620_930# 0.08218f
C130 a_3434_351# a_3567_n217# 0.22378f
C131 a_656_351# a_620_930# 0.24146f
C132 VPWR a_4776_351# 1.11414f
C133 a_750_351# a_656_351# 0.42803f
C134 a_7397_n2523# a_6118_351# 0.11621f
C135 a_745_n2395# a_2026_n1958# 0.23834f
C136 a_2087_n2395# a_620_930# 0.05403f
C137 a_2092_351# a_620_930# 0.04f
C138 VPWR a_4771_n2395# 0.98193f
C139 a_3429_n2395# a_4771_n2395# 0.7336f
C140 a_750_351# a_2092_351# 0.77984f
R0 vctl.n22 vctl.n0 33.8794
R1 vctl.n21 vctl.n20 33.5376
R2 vctl.n6 vctl.n4 24.4981
R3 vctl.n10 vctl.n9 24.4978
R4 vctl.n14 vctl.n13 24.4978
R5 vctl.n18 vctl.n17 24.495
R6 vctl.n6 vctl.n5 24.4894
R7 vctl.n10 vctl.n8 24.488
R8 vctl.n18 vctl.n16 24.4838
R9 vctl.n14 vctl.n12 24.4796
R10 vctl.n3 vctl.n1 24.4574
R11 vctl.n3 vctl.n2 24.4469
R12 vctl.n7 vctl.n3 10.719
R13 vctl.n19 vctl.n18 9.0005
R14 vctl.n15 vctl.n14 9.0005
R15 vctl.n11 vctl.n10 9.0005
R16 vctl.n7 vctl.n6 9.0005
R17 vctl.n21 vctl.n19 1.69764
R18 vctl.n19 vctl.n15 1.68884
R19 vctl.n15 vctl.n11 1.68004
R20 vctl.n11 vctl.n7 1.66496
R21 vctl vctl.n22 0.698214
R22 vctl.n22 vctl.n21 0.569986
R23 VGND.n110 VGND.n36 795000
R24 VGND.n108 VGND.n102 408611
R25 VGND.n178 VGND.n177 36759.9
R26 VGND.n92 VGND.n91 27000
R27 VGND.n91 VGND.n12 27000
R28 VGND.n46 VGND.n12 27000
R29 VGND.n105 VGND.n10 24089.8
R30 VGND.n107 VGND.n106 24089.8
R31 VGND.n109 VGND.n108 22334.8
R32 VGND.n176 VGND.n175 21736.5
R33 VGND.n109 VGND.n101 21565.7
R34 VGND.n47 VGND.n46 20644.2
R35 VGND.n177 VGND.n9 19846.7
R36 VGND.n178 VGND.n8 14324.5
R37 VGND.n179 VGND.n178 11796.7
R38 VGND.n86 VGND.n46 10432.6
R39 VGND.n176 VGND.n8 6890.98
R40 VGND.n92 VGND.n89 6755.73
R41 VGND.n91 VGND.n88 6755.73
R42 VGND.n91 VGND.n90 6755.73
R43 VGND.n87 VGND.n12 6755.73
R44 VGND.n173 VGND.n12 6755.73
R45 VGND.n105 VGND.n18 6068.7
R46 VGND.n106 VGND.n104 6068.7
R47 VGND.n107 VGND.n27 6068.7
R48 VGND.n103 VGND.n10 6068.7
R49 VGND.n175 VGND.n174 6068.7
R50 VGND.n102 VGND.n101 5388.03
R51 VGND.n94 VGND.n93 5194.39
R52 VGND.n93 VGND.n92 4867.89
R53 VGND.n86 VGND.n85 4042.39
R54 VGND.n110 VGND.n109 3958.31
R55 VGND.n104 VGND.n102 3571.26
R56 VGND.n93 VGND.n88 3126.84
R57 VGND.n111 VGND.n110 3045.98
R58 VGND.n85 VGND.n47 3000
R59 VGND.n103 VGND.n8 2384.11
R60 VGND.n104 VGND.n103 2380.84
R61 VGND.n88 VGND.n87 2371.02
R62 VGND.n87 VGND.n86 2282.62
R63 VGND.n57 VGND.n54 1155.83
R64 VGND.n170 VGND.n13 1155.83
R65 VGND.n152 VGND.n25 1155.83
R66 VGND.n135 VGND.n34 1155.83
R67 VGND.n111 VGND.n101 303.187
R68 VGND.n48 VGND.n6 295.591
R69 VGND.n174 VGND.n11 281.534
R70 VGND.n173 VGND.n172 281.534
R71 VGND.n169 VGND.n18 281.534
R72 VGND.n90 VGND.n22 281.534
R73 VGND.n151 VGND.n27 281.534
R74 VGND.n89 VGND.n31 281.534
R75 VGND.n112 VGND.n40 259.877
R76 VGND.n95 VGND.n94 258.901
R77 VGND.n47 VGND.n9 167.286
R78 VGND.n85 VGND.n84 131.024
R79 VGND.n134 VGND.n36 113.647
R80 VGND.n112 VGND.n111 113.186
R81 VGND.n77 VGND.n9 112.975
R82 VGND.n95 VGND.n36 108.236
R83 VGND.n40 VGND.n36 108.23
R84 VGND.n48 VGND.n5 81.1742
R85 VGND.n180 VGND.n6 76.6484
R86 VGND.n177 VGND.n176 22.5473
R87 VGND.n180 VGND.n179 18.3095
R88 VGND.n106 VGND.n105 17.9646
R89 VGND.n108 VGND.n107 17.9646
R90 VGND.n175 VGND.n10 17.9646
R91 VGND.n76 VGND.n56 17.0607
R92 VGND.n119 VGND.n118 17.0177
R93 VGND.n77 VGND.n76 17.0005
R94 VGND.n79 VGND.n78 17.0005
R95 VGND.n78 VGND.n53 17.0005
R96 VGND.n133 VGND.n38 17.0005
R97 VGND.n150 VGND.n29 17.0005
R98 VGND.n168 VGND.n20 17.0005
R99 VGND.n67 VGND.n66 17.0005
R100 VGND.n132 VGND.n131 9.08291
R101 VGND.n124 VGND.n32 9.08291
R102 VGND.n149 VGND.n148 9.08291
R103 VGND.n141 VGND.n23 9.08291
R104 VGND.n158 VGND.n157 9.08291
R105 VGND.n162 VGND.n16 9.08291
R106 VGND.n65 VGND.n64 9.08291
R107 VGND.n113 VGND.n41 9.08291
R108 VGND.n45 VGND.n44 9.07702
R109 VGND.n3 VGND.n0 9.03039
R110 VGND VGND.n183 9.02847
R111 VGND.n126 VGND.n125 9.0005
R112 VGND.n130 VGND.n123 9.0005
R113 VGND.n143 VGND.n142 9.0005
R114 VGND.n147 VGND.n140 9.0005
R115 VGND.n164 VGND.n163 9.0005
R116 VGND.n160 VGND.n159 9.0005
R117 VGND.n62 VGND.n59 9.0005
R118 VGND.n115 VGND.n114 9.0005
R119 VGND.n117 VGND.n116 9.0005
R120 VGND.n99 VGND.n98 9.0005
R121 VGND.n100 VGND.n43 9.0005
R122 VGND.n72 VGND.n71 9.0005
R123 VGND.n70 VGND.n56 9.0005
R124 VGND.n128 VGND.n127 9.0005
R125 VGND.n145 VGND.n144 9.0005
R126 VGND.n166 VGND.n165 9.0005
R127 VGND.n69 VGND.n53 9.0005
R128 VGND.n129 VGND.n38 9.0005
R129 VGND.n146 VGND.n29 9.0005
R130 VGND.n161 VGND.n20 9.0005
R131 VGND.n68 VGND.n67 9.0005
R132 VGND.n2 VGND.n1 9.0005
R133 VGND.n183 VGND.n182 9.0005
R134 VGND.n57 VGND.n52 8.501
R135 VGND.n84 VGND.n83 8.5005
R136 VGND.n97 VGND.n96 8.4728
R137 VGND.n119 VGND.n42 8.4706
R138 VGND.n66 VGND.n61 8.4706
R139 VGND.n168 VGND.n156 8.4706
R140 VGND.n150 VGND.n139 8.4706
R141 VGND.n133 VGND.n122 8.4706
R142 VGND.n74 VGND.n58 8.4706
R143 VGND.n74 VGND.n73 8.4706
R144 VGND.n96 VGND.n45 5.63627
R145 VGND.n136 VGND.n33 5.63396
R146 VGND.n153 VGND.n24 5.63396
R147 VGND.n171 VGND.n17 5.63396
R148 VGND.n136 VGND.n32 5.63382
R149 VGND.n153 VGND.n23 5.63382
R150 VGND.n171 VGND.n16 5.63382
R151 VGND.n119 VGND.n41 5.63382
R152 VGND.n66 VGND.n65 5.63382
R153 VGND.n168 VGND.n157 5.63382
R154 VGND.n150 VGND.n149 5.63382
R155 VGND.n133 VGND.n132 5.63382
R156 VGND.n162 VGND.n14 5.40173
R157 VGND.n113 VGND.n112 5.39607
R158 VGND.n70 VGND.n55 5.39516
R159 VGND.n141 VGND.n26 5.39516
R160 VGND.n124 VGND.n35 5.39513
R161 VGND.n94 VGND.n44 5.36707
R162 VGND.n64 VGND.n63 5.3654
R163 VGND.n158 VGND.n19 5.3654
R164 VGND.n148 VGND.n28 5.3654
R165 VGND.n131 VGND.n37 5.3654
R166 VGND.n77 VGND.n54 5.16623
R167 VGND.n57 VGND.n11 5.16623
R168 VGND.n172 VGND.n13 5.16623
R169 VGND.n170 VGND.n169 5.16623
R170 VGND.n25 VGND.n22 5.16623
R171 VGND.n152 VGND.n151 5.16623
R172 VGND.n34 VGND.n31 5.16623
R173 VGND.n135 VGND.n134 5.16623
R174 VGND VGND.n0 4.5188
R175 VGND.n75 VGND.n57 4.25119
R176 VGND.n174 VGND.n173 3.8748
R177 VGND.n90 VGND.n18 3.8748
R178 VGND.n89 VGND.n27 3.8748
R179 VGND.n80 VGND.n50 3.57718
R180 VGND.n78 VGND.n77 3.4005
R181 VGND.n84 VGND.n5 3.38905
R182 VGND.n182 VGND.n181 3.12829
R183 VGND.n120 VGND.n119 2.95625
R184 VGND.n171 VGND.n15 2.95625
R185 VGND.n154 VGND.n153 2.95625
R186 VGND.n137 VGND.n136 2.95625
R187 VGND.n133 VGND.n30 2.95617
R188 VGND.n150 VGND.n21 2.95617
R189 VGND.n168 VGND.n167 2.95617
R190 VGND.n66 VGND.n51 2.95617
R191 VGND.n83 VGND.n49 2.9539
R192 VGND.n181 VGND.n5 2.83458
R193 VGND.n57 VGND.n55 2.83383
R194 VGND.n77 VGND.n55 2.83383
R195 VGND.n170 VGND.n14 2.83383
R196 VGND.n172 VGND.n14 2.83383
R197 VGND.n152 VGND.n26 2.83383
R198 VGND.n26 VGND.n22 2.83383
R199 VGND.n135 VGND.n35 2.83383
R200 VGND.n35 VGND.n31 2.83383
R201 VGND.n63 VGND.n11 2.83383
R202 VGND.n63 VGND.n54 2.83383
R203 VGND.n169 VGND.n19 2.83383
R204 VGND.n19 VGND.n13 2.83383
R205 VGND.n151 VGND.n28 2.83383
R206 VGND.n28 VGND.n25 2.83383
R207 VGND.n134 VGND.n37 2.83383
R208 VGND.n37 VGND.n34 2.83383
R209 VGND.n172 VGND.n171 2.83383
R210 VGND.n153 VGND.n22 2.83383
R211 VGND.n136 VGND.n31 2.83383
R212 VGND.n136 VGND.n135 2.83383
R213 VGND.n153 VGND.n152 2.83383
R214 VGND.n171 VGND.n170 2.83383
R215 VGND.n134 VGND.n133 2.83383
R216 VGND.n133 VGND.n34 2.83383
R217 VGND.n151 VGND.n150 2.83383
R218 VGND.n150 VGND.n25 2.83383
R219 VGND.n169 VGND.n168 2.83383
R220 VGND.n168 VGND.n13 2.83383
R221 VGND.n66 VGND.n11 2.83383
R222 VGND.n66 VGND.n54 2.83383
R223 VGND.n181 VGND.n180 2.83383
R224 VGND.n181 VGND.n4 2.80958
R225 VGND.n83 VGND.n82 2.73145
R226 VGND.n82 VGND.n7 2.6007
R227 VGND.n96 VGND.n39 2.48001
R228 VGND.n4 VGND.n3 0.962312
R229 VGND.n179 VGND.n7 0.744593
R230 VGND.n129 VGND.n128 0.3701
R231 VGND.n146 VGND.n145 0.3701
R232 VGND.n165 VGND.n161 0.3701
R233 VGND.n69 VGND.n68 0.3701
R234 VGND.n116 VGND.n100 0.3701
R235 VGND.n182 VGND.n2 0.3555
R236 VGND.n3 VGND.n2 0.353
R237 VGND.n53 VGND.n51 0.323287
R238 VGND.n167 VGND.n166 0.323287
R239 VGND.n144 VGND.n21 0.323287
R240 VGND.n127 VGND.n30 0.323287
R241 VGND.n81 VGND.n49 0.308397
R242 VGND.n118 VGND.n39 0.262968
R243 VGND.n82 VGND.n81 0.224343
R244 VGND.n49 VGND.n4 0.195252
R245 VGND.n131 VGND.n130 0.192746
R246 VGND.n126 VGND.n124 0.192746
R247 VGND.n148 VGND.n147 0.192746
R248 VGND.n143 VGND.n141 0.192746
R249 VGND.n160 VGND.n158 0.192746
R250 VGND.n164 VGND.n162 0.192746
R251 VGND.n64 VGND.n59 0.192746
R252 VGND.n71 VGND.n70 0.192746
R253 VGND.n99 VGND.n44 0.192746
R254 VGND.n115 VGND.n113 0.192746
R255 VGND.n130 VGND.n129 0.191392
R256 VGND.n128 VGND.n126 0.191392
R257 VGND.n147 VGND.n146 0.191392
R258 VGND.n145 VGND.n143 0.191392
R259 VGND.n161 VGND.n160 0.191392
R260 VGND.n165 VGND.n164 0.191392
R261 VGND.n68 VGND.n59 0.191392
R262 VGND.n71 VGND.n69 0.191392
R263 VGND.n100 VGND.n99 0.191392
R264 VGND.n116 VGND.n115 0.191392
R265 VGND.n132 VGND.n123 0.163122
R266 VGND.n149 VGND.n140 0.163122
R267 VGND.n159 VGND.n157 0.163122
R268 VGND.n65 VGND.n62 0.163122
R269 VGND.n114 VGND.n41 0.163122
R270 VGND.n163 VGND.n16 0.163122
R271 VGND.n142 VGND.n23 0.163122
R272 VGND.n125 VGND.n32 0.163122
R273 VGND.n138 VGND.n137 0.158669
R274 VGND.n155 VGND.n154 0.158669
R275 VGND.n60 VGND.n15 0.158669
R276 VGND.n121 VGND.n120 0.158669
R277 VGND.n81 VGND.n80 0.158149
R278 VGND.n125 VGND.n33 0.154735
R279 VGND.n142 VGND.n24 0.154735
R280 VGND.n163 VGND.n17 0.154735
R281 VGND.n98 VGND.n45 0.151468
R282 VGND.n123 VGND.n122 0.123672
R283 VGND.n140 VGND.n139 0.123672
R284 VGND.n159 VGND.n156 0.123672
R285 VGND.n62 VGND.n61 0.123672
R286 VGND.n114 VGND.n42 0.123672
R287 VGND.n73 VGND.n72 0.123672
R288 VGND.n58 VGND.n56 0.123672
R289 VGND.n72 VGND.n58 0.121954
R290 VGND.n117 VGND.n42 0.120235
R291 VGND.n98 VGND.n97 0.114798
R292 VGND.n97 VGND.n43 0.111609
R293 VGND.n122 VGND.n121 0.0927349
R294 VGND.n139 VGND.n138 0.0927349
R295 VGND.n156 VGND.n155 0.0927349
R296 VGND.n61 VGND.n60 0.0927349
R297 VGND.n73 VGND.n53 0.0927349
R298 VGND.n127 VGND.n33 0.06234
R299 VGND.n144 VGND.n24 0.06234
R300 VGND.n166 VGND.n17 0.06234
R301 VGND.n183 VGND.n1 0.0597227
R302 VGND.n120 VGND.n39 0.0487297
R303 VGND.n118 VGND.n117 0.04175
R304 VGND.n118 VGND.n43 0.0403551
R305 VGND.n1 VGND.n0 0.0302293
R306 VGND.n7 VGND.n6 0.0072732
R307 VGND.n167 VGND.n15 0.00274058
R308 VGND.n154 VGND.n21 0.00274058
R309 VGND.n137 VGND.n30 0.00274058
R310 VGND.n79 VGND.n51 0.00194262
R311 VGND.n67 VGND.n53 0.00194262
R312 VGND.n166 VGND.n20 0.00194262
R313 VGND.n144 VGND.n29 0.00194262
R314 VGND.n127 VGND.n38 0.00194262
R315 VGND.n76 VGND.n50 0.00170566
R316 VGND.n76 VGND.n75 0.00162501
R317 VGND.n83 VGND.n48 0.00157929
R318 VGND.n75 VGND.n74 0.00137498
R319 VGND.n96 VGND.n95 0.00135895
R320 VGND.n78 VGND.n50 0.00129432
R321 VGND.n119 VGND.n40 0.00111193
R322 VGND.n78 VGND.n52 0.001
R323 VGND.n74 VGND.n52 0.001
R324 VGND.n80 VGND.n79 0.000860656
R325 VGND.n67 VGND.n60 0.000860656
R326 VGND.n155 VGND.n20 0.000860656
R327 VGND.n138 VGND.n29 0.000860656
R328 VGND.n121 VGND.n38 0.000860656
R329 Vout Vout.n1 20.53
R330 Vout.n1 Vout.n0 0.0188902
C141 vctl VGND 11.2953f
C142 Vout VGND 8.14842f
C143 VPWR VGND 11.1055f
C144 m2_7727_571# VGND 0.04717f $ **FLOATING
C145 a_7397_n2523# VGND 0.05072f $ **FLOATING
C146 a_6051_n2525# VGND 0.04654f $ **FLOATING
C147 a_4709_n2525# VGND 0.0474f $ **FLOATING
C148 a_3367_n2525# VGND 0.04814f $ **FLOATING
C149 a_2025_n2525# VGND 0.04567f $ **FLOATING
C150 a_683_n2525# VGND 0.07408f $ **FLOATING
C151 a_6113_n2395# VGND 4.52843f $ **FLOATING
C152 a_4771_n2395# VGND 4.66244f $ **FLOATING
C153 a_3429_n2395# VGND 4.71205f $ **FLOATING
C154 a_2087_n2395# VGND 5.15226f $ **FLOATING
C155 a_745_n2395# VGND 5.27135f $ **FLOATING
C156 a_7398_n1956# VGND 0.75072f $ **FLOATING
C157 a_6052_n1958# VGND 0.8045f $ **FLOATING
C158 a_4710_n1958# VGND 0.81785f $ **FLOATING
C159 a_3368_n1958# VGND 0.82955f $ **FLOATING
C160 a_2026_n1958# VGND 0.82862f $ **FLOATING
C161 a_684_n1958# VGND 0.83893f $ **FLOATING
C162 a_7198_n376# VGND 0.27582f $ **FLOATING
C163 a_6251_n217# VGND 0.65331f $ **FLOATING
C164 a_4909_n217# VGND 0.67139f $ **FLOATING
C165 a_3567_n217# VGND 0.6715f $ **FLOATING
C166 a_2225_n217# VGND 0.67644f $ **FLOATING
C167 a_883_n217# VGND 0.68389f $ **FLOATING
C168 a_7212_321# VGND 0.26455f $ **FLOATING
C169 a_6118_351# VGND 6.88f $ **FLOATING
C170 a_4776_351# VGND 4.93597f $ **FLOATING
C171 a_3434_351# VGND 4.4055f $ **FLOATING
C172 a_2092_351# VGND 4.40424f $ **FLOATING
C173 a_750_351# VGND 4.67142f $ **FLOATING
C174 a_542_269# VGND 6.17341f $ **FLOATING
C175 a_6024_351# VGND 0.05855f $ **FLOATING
C176 a_4682_351# VGND 0.03844f $ **FLOATING
C177 a_3340_351# VGND 0.04051f $ **FLOATING
C178 a_1998_351# VGND 0.04084f $ **FLOATING
C179 a_656_351# VGND 0.05472f $ **FLOATING
C180 a_620_930# VGND 5.65746f $ **FLOATING
.ends
