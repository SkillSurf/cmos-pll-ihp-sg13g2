** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_dff_tb.sch
**.subckt t2_dff_tb
x1 VDD GND D CLK RST Q QN t2_dff
Vs VDD GND 1.2
* noconn Q
* noconn QN
Vdin D GND dc 0 ac 0 pulse(0, 1.2, 0, 50p, 50p, 2.5n, 5n)
Vclk CLK GND dc 0 ac 0 pulse(0, 1.2, 0, 50p, 50p, 1.25n, 2.5n)
Vrst RST GND dc 0 ac 0 pulse(0, 1.2, 0, 50p, 50p, 8n, 15n)
**** begin user architecture code


.param temp=27
.control
save all
tran 10p 15n
write tran_t2_dff.raw
.endc



.lib cornerMOSlv.lib mos_ff

**** end user architecture code
**.ends

* expanding   symbol:  t2_dff.sym # of pins=7
** sym_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_dff.sym
** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_dff.sch
.subckt t2_dff VDD VSS D CLK RST Q QN
*.iopin VSS
*.ipin D
*.ipin RST
*.opin Q
*.iopin VDD
*.opin QN
*.ipin CLK
x3 VDD net1 QN Q VSS t2_nand2
x4 VDD VSS Q net2 RST QN t2_nand3
x1 VDD VSS net4 net5 RST net1 t2_nand3
x2 VDD VSS net1 net5 net3 net2 t2_nand3
x6 VDD net3 net1 net4 VSS t2_nand2
x5 VDD VSS net2 D RST net3 t2_nand3
x7 VDD CLK net5 VSS t2_inverter
.ends


* expanding   symbol:  t2_nand2.sym # of pins=5
** sym_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand2.sym
** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand2.sch
.subckt t2_nand2 VDD inA inB out VSS
*.iopin VSS
*.ipin inA
*.ipin inB
*.opin out
*.iopin VDD
XM1 out inA VDD VDD sg13_lv_pmos w=0.3u l=0.15u ng=1 m=1
XM2 out inB VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
XM3 out inB net1 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM4 net1 inA VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  t2_nand3.sym # of pins=6
** sym_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand3.sym
** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand3.sch
.subckt t2_nand3 VDD VSS inA inB inC out
*.iopin VSS
*.ipin inA
*.ipin inC
*.opin out
*.iopin VDD
*.ipin inB
XM1 out inB VDD VDD sg13_lv_pmos w=0.3u l=0.15u ng=1 m=1
XM2 out inC VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
XM3 out inC net1 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM4 net1 inB net2 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM5 net2 inA VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM0 out inA VDD VDD sg13_lv_pmos w=0.3u l=0.15u ng=1 m=1
.ends


* expanding   symbol:  t2_inverter.sym # of pins=4
** sym_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_inverter.sym
** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_inverter.sch
.subckt t2_inverter VP A Y VN
*.iopin VP
*.iopin VN
*.ipin A
*.opin Y
XM2 Y A VP VP sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
XM1 Y A VN VN sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
