* Extracted by KLayout with SG13G2 LVS runset on : 10/06/2025 10:29

.SUBCKT t2_tie
M$1 1 3 3 1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u PD=1.34u
M$2 4 5 1 1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u PD=1.34u
M$3 6 3 2 2 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u PD=1.28u
M$4 2 5 5 2 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u PD=1.28u
.ENDS t2_tie
