** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_vco_inverter_tb_pulse.sch
**.subckt t2_vco_inverter_tb_pulse Vout
*.opin Vout
Vin Vin GND PULSE(0 1.2 0 1n 1n 10n 20n)
Vdd Vdd GND 1.2
x1 Vdd Vdd Vin Vout GND GND t2_vco_inverter
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt



.param temp=27
.tran 0.1n 100n
.save all


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_vco_inverter.sym # of pins=6
** sym_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_vco_inverter.sym
** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_vco_inverter.sch
.subckt t2_vco_inverter VPWR VPB A Y VNB VGND
*.iopin VPWR
*.iopin VGND
*.ipin A
*.opin Y
*.iopin VPB
*.iopin VNB
XM2 Y A VPWR VPB sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
XM1 Y A VGND VNB sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
