* Extracted by KLayout with SG13G2 LVS runset on : 13/06/2025 02:42

.SUBCKT t2_bias
M$1 2 4 6 1 sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=4.3u PD=4.3u
M$6 2 4 4 1 sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=4.3u PD=4.3u
M$11 2 4 10 1 sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=4.3u PD=4.3u
M$16 2 3 4 1 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
M$17 6 10 7 1 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.095p PS=1.68u PD=0.88u
M$18 7 5 8 1 sg13_lv_nmos L=0.15u W=0.5u AS=0.095p AD=0.17p PS=0.88u PD=1.68u
M$19 10 10 12 9 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.095p PS=1.68u PD=0.88u
M$20 12 12 14 9 sg13_lv_pmos L=0.15u W=0.5u AS=0.095p AD=0.17p PS=0.88u PD=1.68u
M$21 10 13 14 9 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
M$22 6 15 14 9 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
M$23 14 6 6 9 sg13_lv_pmos L=1u W=1u AS=0.34p AD=0.34p PS=4.3u PD=4.3u
M$28 11 6 4 9 sg13_lv_pmos L=1u W=1u AS=0.34p AD=0.34p PS=4.3u PD=4.3u
R$33 11 14 rhigh w=0.5u l=0.5u ps=0 b=0 m=1
.ENDS t2_bias
