* Extracted by KLayout with SG13G2 LVS runset on : 18/07/2025 17:08

.SUBCKT t2_pmos$1
.ENDS t2_pmos$1

.SUBCKT t2_nmos$1
.ENDS t2_nmos$1

.SUBCKT pmos_bulk$1
.ENDS pmos_bulk$1

.SUBCKT 11Stage_vco_new
X$1 1 15 1 cmim$1
X$2 2 1 35 15 15 1 35 15 35 15 2 t2_inverter_buffer$1
X$3 1 11 1 cmim$1
X$4 1 14 1 cmim$1
X$5 1 34 1 cmim$1
X$6 1 16 1 cmim$1
X$7 1 35 1 cmim$1
X$8 1 12 1 cmim$1
X$9 1 35 1 cmim$1
X$10 1 13 1 cmim$1
X$11 1 31 1 cmim$1
X$12 1 9 1 cmim$1
X$13 1 32 1 cmim$1
X$14 1 33 1 cmim$1
X$15 1 22 1 25 nmos$3$2
X$16 22 1 1 25 nmos$3$2
X$17 20 1 1 25 nmos$6
X$18 21 1 1 25 nmos$6
X$19 19 1 1 25 nmos$6
X$20 18 1 1 25 nmos$6
X$21 17 1 1 25 nmos$6
X$22 10 1 1 25 nmos$6
X$23 30 1 1 25 nmos$6
X$24 29 1 1 25 nmos$6
X$25 27 1 1 25 nmos$6
X$26 1 17 1 25 nmos$6
X$27 1 18 1 25 nmos$6
X$28 1 20 1 25 nmos$6
X$29 1 19 1 25 nmos$6
X$30 1 10 1 25 nmos$6
X$31 1 26 1 25 nmos$6
X$32 1 28 1 25 nmos$6
X$33 1 30 1 25 nmos$6
X$34 1 29 1 25 nmos$6
X$35 1 27 1 25 nmos$6
X$36 1 21 1 25 nmos$6
X$37 26 1 1 25 nmos$6
X$38 28 1 1 25 nmos$6
X$39 2 8 10 2 1 pmos$3$1
X$40 8 2 10 2 1 pmos$3$1
X$41 2 8 10 2 1 pmos$3$1
X$42 8 2 10 2 1 pmos$3$1
X$43 2 10 10 2 1 pmos$6
X$44 10 2 10 2 1 pmos$6
X$45 2 10 10 2 1 pmos$6
X$46 10 2 10 2 1 pmos$6
X$47 5 2 10 2 1 pmos$6
X$48 2 5 10 2 1 pmos$6
X$49 2 5 10 2 1 pmos$6
X$50 5 2 10 2 1 pmos$6
X$51 3 2 10 2 1 pmos$6
X$52 2 3 10 2 1 pmos$6
X$53 2 3 10 2 1 pmos$6
X$54 3 2 10 2 1 pmos$6
X$55 4 2 10 2 1 pmos$6
X$56 2 4 10 2 1 pmos$6
X$57 2 4 10 2 1 pmos$6
X$58 4 2 10 2 1 pmos$6
X$59 6 2 10 2 1 pmos$6
X$60 2 6 10 2 1 pmos$6
X$61 2 6 10 2 1 pmos$6
X$62 6 2 10 2 1 pmos$6
X$63 7 2 10 2 1 pmos$6
X$64 2 7 10 2 1 pmos$6
X$65 2 7 10 2 1 pmos$6
X$66 7 2 10 2 1 pmos$6
X$67 38 2 10 2 1 pmos$6
X$68 2 38 10 2 1 pmos$6
X$69 2 38 10 2 1 pmos$6
X$70 38 2 10 2 1 pmos$6
X$71 36 2 10 2 1 pmos$6
X$72 2 36 10 2 1 pmos$6
X$73 2 36 10 2 1 pmos$6
X$74 36 2 10 2 1 pmos$6
X$75 37 2 10 2 1 pmos$6
X$76 2 37 10 2 1 pmos$6
X$77 2 37 10 2 1 pmos$6
X$78 37 2 10 2 1 pmos$6
X$79 39 2 10 2 1 pmos$6
X$80 2 39 10 2 1 pmos$6
X$81 2 39 10 2 1 pmos$6
X$82 39 2 10 2 1 pmos$6
X$83 40 2 10 2 1 pmos$6
X$84 2 40 10 2 1 pmos$6
X$85 2 40 10 2 1 pmos$6
X$86 40 2 10 2 1 pmos$6
X$87 1 36 2 31 16 28 VCO_1$1
X$88 17 16 1 11 nmos$2$2
X$89 16 17 1 11 nmos$2$2
X$90 1 37 2 32 31 29 VCO_1$1
X$91 18 11 1 12 nmos$2$2
X$92 11 18 1 12 nmos$2$2
X$93 1 38 2 33 32 30 VCO_1$1
X$94 19 12 1 13 nmos$2$2
X$95 12 19 1 13 nmos$2$2
X$96 1 39 2 34 33 26 VCO_1$1
X$97 20 13 1 14 nmos$2$2
X$98 13 20 1 14 nmos$2$2
X$99 1 40 2 15 34 27 VCO_1$1
X$100 21 14 1 9 nmos$2$2
X$101 14 21 1 9 nmos$2$2
X$102 9 22 1 15 nmos$2$2
X$103 22 9 1 15 nmos$2$2
X$104 9 8 15 2 1 pmos$2$2
X$105 8 9 15 2 1 pmos$2$2
X$106 8 9 15 2 1 pmos$2$2
X$107 9 8 15 2 1 pmos$2$2
X$108 14 7 9 2 1 pmos$2$2
X$109 7 14 9 2 1 pmos$2$2
X$110 7 14 9 2 1 pmos$2$2
X$111 14 7 9 2 1 pmos$2$2
X$112 13 6 14 2 1 pmos$2$2
X$113 6 13 14 2 1 pmos$2$2
X$114 6 13 14 2 1 pmos$2$2
X$115 13 6 14 2 1 pmos$2$2
X$116 11 4 12 2 1 pmos$2$2
X$117 4 11 12 2 1 pmos$2$2
X$118 4 11 12 2 1 pmos$2$2
X$119 11 4 12 2 1 pmos$2$2
X$120 16 3 11 2 1 pmos$2$2
X$121 3 16 11 2 1 pmos$2$2
X$122 3 16 11 2 1 pmos$2$2
X$123 16 3 11 2 1 pmos$2$2
X$124 12 5 13 2 1 pmos$2$2
X$125 5 12 13 2 1 pmos$2$2
X$126 5 12 13 2 1 pmos$2$2
X$127 12 5 13 2 1 pmos$2$2
M$1 1 25 27 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p PS=1.28u PD=0.74u
M$2 27 25 1 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p PS=0.74u PD=1.28u
M$3 1 25 26 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p PS=1.28u PD=0.74u
M$4 26 25 1 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p PS=0.74u PD=1.28u
M$5 1 25 30 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p PS=1.28u PD=0.74u
M$6 30 25 1 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p PS=0.74u PD=1.28u
M$7 1 25 29 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p PS=1.28u PD=0.74u
M$8 29 25 1 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p PS=0.74u PD=1.28u
M$9 1 25 28 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p PS=1.28u PD=0.74u
M$10 28 25 1 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p PS=0.74u PD=1.28u
M$11 1 25 22 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p PS=1.28u PD=0.74u
M$12 22 25 1 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p PS=0.74u PD=1.28u
M$13 1 25 21 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p PS=1.28u PD=0.74u
M$14 21 25 1 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p PS=0.74u PD=1.28u
M$15 1 25 20 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p PS=1.28u PD=0.74u
M$16 20 25 1 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p PS=0.74u PD=1.28u
M$17 1 25 19 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p PS=1.28u PD=0.74u
M$18 19 25 1 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p PS=0.74u PD=1.28u
M$19 20 14 13 1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p PS=1.34u
+ PD=0.74u
M$20 13 14 20 1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p PS=0.74u
+ PD=1.34u
M$21 1 25 10 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p PS=1.28u PD=0.74u
M$22 10 25 1 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p PS=0.74u PD=1.28u
M$23 19 13 12 1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p PS=1.34u
+ PD=0.74u
M$24 12 13 19 1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p PS=0.74u
+ PD=1.34u
M$25 18 12 11 1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p PS=1.34u
+ PD=0.74u
M$26 11 12 18 1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p PS=0.74u
+ PD=1.34u
M$27 17 11 16 1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p PS=1.34u
+ PD=0.74u
M$28 16 11 17 1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p PS=0.74u
+ PD=1.34u
M$29 22 15 9 1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p PS=1.34u
+ PD=0.74u
M$30 9 15 22 1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p PS=0.74u
+ PD=1.34u
M$31 21 9 14 1 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p PS=1.34u
+ PD=0.74u
M$32 14 9 21 1 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p PS=0.74u
+ PD=1.34u
M$33 1 25 18 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p PS=1.28u PD=0.74u
M$34 18 25 1 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p PS=0.74u PD=1.28u
M$35 1 25 17 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.066p PS=1.28u PD=0.74u
M$36 17 25 1 1 sg13_lv_nmos L=0.13u W=0.3u AS=0.066p AD=0.102p PS=0.74u PD=1.28u
M$37 37 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p PS=0.745u
+ PD=0.74u
M$38 2 10 37 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$39 37 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.104p PS=0.74u PD=1.34u
M$40 37 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p PS=0.745u
+ PD=1.34u
M$41 36 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p PS=0.745u
+ PD=0.74u
M$42 2 10 36 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$43 36 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.104p PS=0.74u PD=1.34u
M$44 36 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p PS=0.745u
+ PD=1.34u
M$45 40 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p PS=0.745u
+ PD=0.74u
M$46 2 10 40 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$47 40 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.104p PS=0.74u PD=1.34u
M$48 40 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p PS=0.745u
+ PD=1.34u
M$49 39 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p PS=0.745u
+ PD=0.74u
M$50 2 10 39 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$51 39 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.104p PS=0.74u PD=1.34u
M$52 39 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p PS=0.745u
+ PD=1.34u
M$53 9 15 8 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.1075p PS=0.745u
+ PD=1.34u
M$54 8 15 9 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p PS=1.34u
+ PD=0.74u
M$55 9 15 8 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.0625p PS=0.74u
+ PD=0.74u
M$56 9 15 8 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.0625p PS=0.745u
+ PD=0.74u
M$57 14 9 7 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.1075p PS=0.745u
+ PD=1.34u
M$58 7 9 14 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p PS=1.34u
+ PD=0.74u
M$59 14 9 7 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.0625p PS=0.74u
+ PD=0.74u
M$60 14 9 7 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.0625p PS=0.745u
+ PD=0.74u
M$61 8 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p PS=0.745u
+ PD=1.34u
M$62 2 10 8 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.104p AD=0.059p PS=1.34u PD=0.74u
M$63 8 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$64 8 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p PS=0.745u
+ PD=0.74u
M$65 6 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p PS=0.745u
+ PD=1.34u
M$66 2 10 6 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.104p AD=0.059p PS=1.34u PD=0.74u
M$67 6 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$68 6 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p PS=0.745u
+ PD=0.74u
M$69 7 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p PS=0.745u
+ PD=1.34u
M$70 2 10 7 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.104p AD=0.059p PS=1.34u PD=0.74u
M$71 7 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$72 7 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p PS=0.745u
+ PD=0.74u
M$73 2 10 10 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.104p AD=0.059p PS=1.34u PD=0.74u
M$74 10 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$75 2 10 10 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.05975p PS=0.74u
+ PD=0.745u
M$76 10 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p PS=0.745u
+ PD=1.34u
M$77 12 13 5 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.1075p PS=0.745u
+ PD=1.34u
M$78 5 13 12 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p PS=1.34u
+ PD=0.74u
M$79 12 13 5 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.0625p PS=0.74u
+ PD=0.74u
M$80 12 13 5 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.0625p PS=0.745u
+ PD=0.74u
M$81 38 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p PS=0.745u
+ PD=0.74u
M$82 2 10 38 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$83 38 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.104p PS=0.74u PD=1.34u
M$84 38 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p PS=0.745u
+ PD=1.34u
M$85 11 12 4 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.1075p PS=0.745u
+ PD=1.34u
M$86 4 12 11 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p PS=1.34u
+ PD=0.74u
M$87 11 12 4 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.0625p PS=0.74u
+ PD=0.74u
M$88 11 12 4 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.0625p PS=0.745u
+ PD=0.74u
M$89 5 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p PS=0.745u
+ PD=1.34u
M$90 2 10 5 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.104p AD=0.059p PS=1.34u PD=0.74u
M$91 5 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$92 5 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p PS=0.745u
+ PD=0.74u
M$93 3 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p PS=0.745u
+ PD=1.34u
M$94 2 10 3 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.104p AD=0.059p PS=1.34u PD=0.74u
M$95 3 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$96 3 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p PS=0.745u
+ PD=0.74u
M$97 4 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.104p PS=0.745u
+ PD=1.34u
M$98 2 10 4 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.104p AD=0.059p PS=1.34u PD=0.74u
M$99 4 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$100 4 10 2 2 sg13_lv_pmos L=0.13u W=0.2u AS=0.05975p AD=0.059p PS=0.745u
+ PD=0.74u
M$101 13 14 6 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.1075p PS=0.745u
+ PD=1.34u
M$102 6 14 13 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p PS=1.34u
+ PD=0.74u
M$103 13 14 6 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.0625p PS=0.74u
+ PD=0.74u
M$104 13 14 6 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.0625p PS=0.745u
+ PD=0.74u
M$105 16 11 3 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.1075p PS=0.745u
+ PD=1.34u
M$106 3 11 16 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p PS=1.34u
+ PD=0.74u
M$107 16 11 3 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.0625p PS=0.74u
+ PD=0.74u
M$108 16 11 3 2 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.0625p PS=0.745u
+ PD=0.74u
.ENDS 11Stage_vco_new

.SUBCKT nmos$3$2 1 2 3 4
.ENDS nmos$3$2

.SUBCKT pmos$3$1 1 2 3 4 5
.ENDS pmos$3$1

.SUBCKT t2_inverter_buffer$1 1 2 3 4 5 6 7 8 9 10 11
X$1 7 1 5 11 6 pmos$6
X$2 1 9 5 11 6 pmos$6
X$3 1 7 5 11 6 pmos$6
X$4 9 1 5 11 6 pmos$6
X$5 3 2 6 4 nmos$2$2
X$6 2 3 6 4 nmos$2$2
M$1 2 4 3 6 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p PS=1.34u PD=0.74u
M$2 3 4 2 6 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p PS=0.74u PD=1.34u
M$3 1 5 9 11 sg13_lv_pmos L=0.13u W=0.2u AS=0.104p AD=0.059p PS=1.34u PD=0.74u
M$4 9 5 1 11 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$5 1 5 7 11 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.059p PS=0.74u PD=0.74u
M$6 7 5 1 11 sg13_lv_pmos L=0.13u W=0.2u AS=0.059p AD=0.104p PS=0.74u PD=1.34u
.ENDS t2_inverter_buffer$1

.SUBCKT nmos$6 1 2 3 4
.ENDS nmos$6

.SUBCKT cmim$1 1 2 3
C$1 3 2 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
.ENDS cmim$1

.SUBCKT VCO_1$1 1 2 3 4 5 6
X$1 3 1 4 5 6 2 T2_Inverter$1
X$2 1 6 nmos_bulk$1
.ENDS VCO_1$1

.SUBCKT pmos$6 1 2 3 4 5
.ENDS pmos$6

.SUBCKT nmos_bulk$1 1 2
.ENDS nmos_bulk$1

.SUBCKT T2_Inverter$1 1 2 3 4 5 6
X$1 6 3 4 1 2 pmos$2$2
X$2 3 6 4 1 2 pmos$2$2
X$3 3 6 4 1 2 pmos$2$2
X$4 6 3 4 1 2 pmos$2$2
X$5 5 3 2 4 nmos$2$2
X$6 3 5 2 4 nmos$2$2
M$1 5 4 3 2 sg13_lv_nmos L=0.13u W=0.25u AS=0.1075p AD=0.0625p PS=1.34u PD=0.74u
M$2 3 4 5 2 sg13_lv_nmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p PS=0.74u PD=1.34u
M$3 3 4 6 1 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.0625p PS=0.745u
+ PD=0.74u
M$4 6 4 3 1 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.0625p PS=0.74u PD=0.74u
M$5 3 4 6 1 sg13_lv_pmos L=0.13u W=0.25u AS=0.0625p AD=0.1075p PS=0.74u PD=1.34u
M$6 3 4 6 1 sg13_lv_pmos L=0.13u W=0.25u AS=0.06325p AD=0.1075p PS=0.745u
+ PD=1.34u
.ENDS T2_Inverter$1

.SUBCKT nmos$2$2 1 2 3 4
.ENDS nmos$2$2

.SUBCKT pmos$2$2 1 2 3 4 5
.ENDS pmos$2$2
