* Extracted by KLayout with SG13G2 LVS runset on : 10/06/2025 18:09

.SUBCKT t2_or2
M$1 3 4 5 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u PD=0.74u
M$2 5 4 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u PD=1.34u
M$3 6 3 7 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u PD=0.74u
M$4 7 8 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u PD=1.34u
M$5 8 9 10 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$6 10 9 2 2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$7 1 4 3 1 sg13_lv_pmos L=0.13u W=0.6u AS=0.159p AD=0.159p PS=1.96u PD=1.96u
M$9 1 3 6 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$10 6 8 1 1 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$11 1 9 8 1 sg13_lv_pmos L=0.13u W=0.6u AS=0.159p AD=0.159p PS=1.96u PD=1.96u
.ENDS t2_or2
