** sch_path: /foss/designs/Team2/3NAND/3NAND_tb.sch
**.subckt 3NAND_tb Vout
*.opin Vout
Vin VB GND dc 0 ac 0 pulse(0, 1.2, 0, 100p, 100p, 8n, 16n)
Vin1 VA GND dc 0 ac 0 pulse(0, 1.2, 2n, 100p, 100p, 2n, 4n)
C1 Vout GND 100f m=1
x1 Vout VA VB VC 3NAND
Vin2 VC GND dc 0 ac 0 pulse(0, 1.2, 5n, 0.8n, 0.8n, 5n, 10n)
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt



.param temp=27
.control
save all
tran 50p 20n
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/Team2/3NAND/3NAND.sym # of pins=4
** sym_path: /foss/designs/Team2/3NAND/3NAND.sym
** sch_path: /foss/designs/Team2/3NAND/3NAND.sch
.subckt 3NAND Y A B C
*.ipin A
*.ipin B
*.ipin C
*.opin Y
XM1 Y A Vdd Vdd sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM2 Y B Vdd Vdd sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM3 Y C Vdd Vdd sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM4 Y A net1 GND sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM5 net1 B net2 GND sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM6 net2 C GND GND sg13_lv_nmos w=1u l=0.13u ng=1 m=1
V1 Vdd GND 1.2
.ends

.GLOBAL GND
.end
