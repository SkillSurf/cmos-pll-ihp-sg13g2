** sch_path: /foss/designs/iic-osic-tools/cmos-pll-ihp-sg13g2/Combined_Design/design_data/xschem/charge_pump_wo_lpf_tb.sch
**.subckt charge_pump_wo_lpf_tb
V1 VDD GND 1.2
V4 up GND PULSE(0 1.2 .2NS .2NS .2NS 0.02NS 10NS)
V5 down GND PULSE(0 1.2 .2NS .2NS .2NS 2NS 10NS)
x2 VDD bias_p up vout_cp down bias_n GND charge_pump
x3 VDD VDD GND GND net1 bias_n bias_p net2 Bias_gen
V7 net1 GND 1.2
V8 net2 GND 0
C1 vout_cp GND 100f ic=0.5 m=1
**** begin user architecture code


.param temp=27
.tran 1n 100n uic
.save all


 .lib cornerMOSlv.lib mos_tt


.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ_stat

**** end user architecture code
**.ends

* expanding   symbol:  charge_pump.sym # of pins=7
** sym_path: /foss/designs/iic-osic-tools/cmos-pll-ihp-sg13g2/Combined_Design/design_data/xschem/charge_pump.sym
** sch_path: /foss/designs/iic-osic-tools/cmos-pll-ihp-sg13g2/Combined_Design/design_data/xschem/charge_pump.sch
.subckt charge_pump VP bias_p up vout down bias_n VN
*.ipin bias_p
*.ipin up
*.ipin down
*.ipin bias_n
*.iopin VN
*.iopin VP
*.opin vout
XM1 net1 bias_n VN VN sg13_lv_nmos w=1.2u l=0.13u ng=1 m=1
XM2 vout down net1 VN sg13_lv_nmos w=1.2u l=0.13u ng=1 m=1
XM3 vout net3 net2 VP sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM4 net2 bias_p VP VP sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
x1 VP up net3 VN inverter
.ends


* expanding   symbol:  Bias_gen.sym # of pins=8
** sym_path: /foss/designs/iic-osic-tools/cmos-pll-ihp-sg13g2/Combined_Design/design_data/xschem/Bias_gen.sym
** sch_path: /foss/designs/iic-osic-tools/cmos-pll-ihp-sg13g2/Combined_Design/design_data/xschem/Bias_gen.sch
.subckt Bias_gen VPWR VPB VGND VNB en bias_n bias_p enb
*.ipin en
*.opin bias_n
*.iopin VNB
*.iopin VGND
*.iopin VPB
*.iopin VPWR
*.ipin enb
*.opin bias_p
XM1 bias_p kick kick_sw VNB sg13_lv_nmos w=0.5u l=0.15u ng=1 m=1
XM2 kick_sw en VGND VNB sg13_lv_nmos w=0.5u l=0.15u ng=1 m=1
XM3 kick bias_n VGND VNB sg13_lv_nmos w=1.0u l=1.0u ng=1 m=1
XM4 bias_p bias_n net1 VNB sg13_lv_nmos w=1.0u l=1.0u ng=1 m=1
XM5 bias_n enb VGND VNB sg13_lv_nmos w=0.5u l=0.15u ng=1 m=1
XM6 bias_n bias_n VGND VNB sg13_lv_nmos w=1.0u l=1.0u ng=1 m=1
XM7 kick kick dio_mid VPB sg13_lv_pmos w=0.5u l=0.15u ng=1 m=1
XM8 bias_p bias_p VPWR VPB sg13_lv_pmos w=2.0u l=1.0u ng=1 m=1
XM9 bias_p en VPWR VPB sg13_lv_pmos w=0.5u l=0.15u ng=1 m=1
XM10 bias_n bias_p res_bot VPB sg13_lv_pmos w=4.0u l=1.0u ng=1 m=1
XM11 kick en VPWR VPB sg13_lv_pmos w=0.5u l=0.15u ng=1 m=1
XM12 dio_mid dio_mid VPWR VPB sg13_lv_pmos w=0.5u l=0.15u ng=1 m=1
XR1 res_bot VPWR sub! rhigh w=1.0e-6 l=12.0e-6 m=1 b=0
XR2 VGND net1 sub! rhigh w=1.0e-6 l=12.0e-6 m=1 b=0
.ends


* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /foss/designs/iic-osic-tools/cmos-pll-ihp-sg13g2/Combined_Design/design_data/xschem/inverter.sym
** sch_path: /foss/designs/iic-osic-tools/cmos-pll-ihp-sg13g2/Combined_Design/design_data/xschem/inverter.sch
.subckt inverter VP IN OUT VN
*.iopin VN
*.iopin VP
*.ipin IN
*.opin OUT
XM1 OUT IN VN VN sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM2 OUT IN VP VP sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
