** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_charge_pump.sch
.subckt t2_charge_pump VPWR VPB VGND VNB out up down bias_p bias_n
*.PININFO VPWR:B up:I out:O VPB:B VGND:B VNB:B down:I bias_p:I bias_n:I
M1 i_down bias_n VGND VNB sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
M2 out down i_down VNB sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M3 i_up bias_p VPWR VPB sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
M4 out net1 i_up VPB sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
x1 VPWR up net1 VGND t2_inverter
.ends

* expanding   symbol:  t2_inverter.sym # of pins=4
** sym_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_inverter.sym
** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_inverter.sch
.subckt t2_inverter VP A Y VN
*.PININFO VP:B VN:B A:I Y:O
M2 Y A VP VP sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M1 Y A VN VN sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends

