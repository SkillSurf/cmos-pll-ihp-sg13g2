** sch_path: /foss/designs/t2_PFD/t2_PFD_tb.sch
**.subckt t2_PFD_tb
x1 vdd up GND down ref_clk vco_clk t2_PFD
V1 vdd GND 1.2
V2 ref_clk GND PULSE(0 1.2 0 50p 50p 2.5n 5n
V3 vco_clk GND PULSE(0 1.2 1n 50p 50p 2.5n 5n
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt



.param temp=27
.control
save all
tran 10p 40n
write tran_pfd_t2.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  t2_PFD.sym # of pins=6
** sym_path: /foss/designs/t2_PFD/t2_PFD.sym
** sch_path: /foss/designs/t2_PFD/t2_PFD.sch
.subckt t2_PFD vdd up vss down ref_clk vco_clk
*.iopin vdd
*.ipin ref_clk
*.iopin vss
*.ipin vco_clk
*.opin up
*.opin down
XM1 net2 vco_clk vss vss sg13_lv_nmos w=0.36u l=0.15u ng=1 m=1
XM4 net1 ref_clk net2 vss sg13_lv_nmos w=1.8u l=0.15u ng=1 m=1
XM5 net3 ref_clk net1 vss sg13_lv_nmos w=0.84u l=0.15u ng=1 m=1
XM9 net3 ref_clk ref_clk vdd sg13_lv_pmos w=0.64u l=0.15u ng=1 m=1
XM11 net7 net3 vss vss sg13_lv_nmos w=0.36u l=0.15u ng=1 m=1
XM12 vdd net3 net7 vdd sg13_lv_pmos w=0.72u l=0.15u ng=1 m=1
XM13 up net7 vss vss sg13_lv_nmos w=0.48u l=0.15u ng=1 m=1
XM14 vdd net7 up vdd sg13_lv_pmos w=0.96u l=0.15u ng=1 m=1
XM3 net1 ref_clk vdd vdd sg13_lv_pmos w=0.64u l=0.15u ng=1 m=1
XM6 net4 vco_clk vdd vdd sg13_lv_pmos w=0.64u l=0.15u ng=1 m=1
XM7 net4 vco_clk net5 vss sg13_lv_nmos w=1.8u l=0.15u ng=1 m=1
XM19 net5 ref_clk vss vss sg13_lv_nmos w=0.36u l=0.15u ng=1 m=1
XM8 net6 vco_clk net4 vss sg13_lv_nmos w=0.84u l=0.15u ng=1 m=1
XM10 net6 vco_clk vco_clk vdd sg13_lv_pmos w=0.64u l=0.15u ng=1 m=1
XM15 vdd net6 net8 vdd sg13_lv_pmos w=0.72u l=0.15u ng=1 m=1
XM16 net8 net6 vss vss sg13_lv_nmos w=0.36u l=0.15u ng=1 m=1
XM17 vdd net8 down vdd sg13_lv_pmos w=0.96u l=0.15u ng=1 m=1
XM18 down net8 vss vss sg13_lv_nmos w=0.48u l=0.15u ng=1 m=1
.ends

.GLOBAL GND
.end
