** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_dff.sch
.subckt t2_dff VDD VSS D CLK RST Q QN
*.PININFO VSS:B D:I RST:I Q:O VDD:B QN:O CLK:I
x3 VDD net1 QN Q VSS t2_nand2
x4 VDD VSS Q net2 RST QN t2_nand3
x1 VDD VSS net4 net5 RST net1 t2_nand3
x2 VDD VSS net1 net5 net3 net2 t2_nand3
x6 VDD net3 net1 net4 VSS t2_nand2
x5 VDD VSS net2 D RST net3 t2_nand3
x7 VDD CLK net5 VSS t2_inverter
.ends

* expanding   symbol:  t2_nand2.sym # of pins=5
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand2.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand2.sch
.subckt t2_nand2 VDD inA inB out VSS
*.PININFO VSS:B inA:I inB:I out:O VDD:B
M1 out inA VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M2 out inB VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M3 out inB net1 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M4 net1 inA VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  t2_nand3.sym # of pins=6
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand3.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand3.sch
.subckt t2_nand3 VDD VSS inA inB inC out
*.PININFO VSS:B inA:I inC:I out:O VDD:B inB:I
M1 out inB VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M2 out inC VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M3 out inC net1 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M4 net1 inB net2 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M5 net2 inA VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M0 out inA VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  t2_inverter.sym # of pins=4
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_inverter.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_inverter.sch
.subckt t2_inverter VP A Y VN
*.PININFO VP:B VN:B A:I Y:O
M2 Y A VP VP sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M1 Y A VN VN sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends

