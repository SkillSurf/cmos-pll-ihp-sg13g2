* Extracted by KLayout with SG13G2 LVS runset on : 10/06/2025 13:15

.SUBCKT VCO
M$1 \$1 \$3 \$4 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$2 \$4 \$3 \$1 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p PS=0.74u
+ PD=0.74u
M$3 \$1 \$3 \$4 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p PS=0.74u
+ PD=0.74u
M$4 \$4 \$3 \$1 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$5 \$1 \$3 \$5 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$6 \$5 \$3 \$1 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p PS=0.74u
+ PD=0.74u
M$7 \$1 \$3 \$5 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p PS=0.74u
+ PD=0.74u
M$8 \$5 \$3 \$1 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$9 \$1 \$3 \$6 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$10 \$6 \$3 \$1 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p
+ PS=0.74u PD=0.74u
M$11 \$1 \$3 \$6 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p
+ PS=0.74u PD=0.74u
M$12 \$6 \$3 \$1 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p
+ PS=0.74u PD=1.34u
M$13 \$1 \$3 \$7 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p
+ PS=1.34u PD=0.74u
M$14 \$7 \$3 \$1 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p
+ PS=0.74u PD=0.74u
M$15 \$1 \$3 \$7 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p
+ PS=0.74u PD=0.74u
M$16 \$7 \$3 \$1 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p
+ PS=0.74u PD=1.34u
M$17 \$1 \$3 \$8 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p
+ PS=1.34u PD=0.74u
M$18 \$8 \$3 \$1 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p
+ PS=0.74u PD=0.74u
M$19 \$1 \$3 \$8 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p
+ PS=0.74u PD=0.74u
M$20 \$8 \$3 \$1 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p
+ PS=0.74u PD=1.34u
M$21 \$1 \$3 \$9 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p
+ PS=1.34u PD=0.74u
M$22 \$9 \$3 \$1 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p
+ PS=0.74u PD=0.74u
M$23 \$1 \$3 \$9 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p
+ PS=0.74u PD=0.74u
M$24 \$9 \$3 \$1 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p
+ PS=0.74u PD=1.34u
M$25 \$5 \$2 \$16 \$1 sg13_lv_nmos L=0.13u W=0.155u AS=0.10085p AD=0.05585p
+ PS=1.34u PD=0.74u
M$26 \$16 \$2 \$23 \$1 sg13_lv_nmos L=0.13u W=0.155u AS=0.05585p AD=0.10085p
+ PS=0.74u PD=1.34u
M$27 \$6 \$16 \$17 \$1 sg13_lv_nmos L=0.13u W=0.155u AS=0.10085p AD=0.05585p
+ PS=1.34u PD=0.74u
M$28 \$17 \$16 \$25 \$1 sg13_lv_nmos L=0.13u W=0.155u AS=0.05585p AD=0.10085p
+ PS=0.74u PD=1.34u
M$29 \$7 \$17 \$18 \$1 sg13_lv_nmos L=0.13u W=0.155u AS=0.10085p AD=0.05585p
+ PS=1.34u PD=0.74u
M$30 \$18 \$17 \$29 \$1 sg13_lv_nmos L=0.13u W=0.155u AS=0.05585p AD=0.10085p
+ PS=0.74u PD=1.34u
M$31 \$8 \$18 \$19 \$1 sg13_lv_nmos L=0.13u W=0.155u AS=0.10085p AD=0.05585p
+ PS=1.34u PD=0.74u
M$32 \$19 \$18 \$32 \$1 sg13_lv_nmos L=0.13u W=0.155u AS=0.05585p AD=0.10085p
+ PS=0.74u PD=1.34u
M$33 \$9 \$19 \$20 \$1 sg13_lv_nmos L=0.13u W=0.155u AS=0.10085p AD=0.05585p
+ PS=1.34u PD=0.74u
M$34 \$20 \$19 \$28 \$1 sg13_lv_nmos L=0.13u W=0.155u AS=0.05585p AD=0.10085p
+ PS=0.74u PD=1.34u
M$35 \$1 \$20 \$2 \$1 sg13_lv_nmos L=0.13u W=0.155u AS=0.10085p AD=0.05585p
+ PS=1.34u PD=0.74u
M$36 \$2 \$20 \$21 \$1 sg13_lv_nmos L=0.13u W=0.155u AS=0.05585p AD=0.10085p
+ PS=0.74u PD=1.34u
M$37 \$33 \$2 \$16 \$45 sg13_lv_pmos L=0.13u W=0.18u AS=0.1026p AD=0.0576p
+ PS=1.34u PD=0.74u
M$38 \$16 \$2 \$33 \$45 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.0576p
+ PS=0.74u PD=0.74u
M$39 \$33 \$2 \$16 \$45 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.0576p
+ PS=0.74u PD=0.74u
M$40 \$16 \$2 \$33 \$45 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.1026p
+ PS=0.74u PD=1.34u
M$41 \$34 \$16 \$17 \$47 sg13_lv_pmos L=0.13u W=0.18u AS=0.1026p AD=0.0576p
+ PS=1.34u PD=0.74u
M$42 \$17 \$16 \$34 \$47 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.0576p
+ PS=0.74u PD=0.74u
M$43 \$34 \$16 \$17 \$47 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.0576p
+ PS=0.74u PD=0.74u
M$44 \$17 \$16 \$34 \$47 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.1026p
+ PS=0.74u PD=1.34u
M$45 \$35 \$17 \$18 \$48 sg13_lv_pmos L=0.13u W=0.18u AS=0.1026p AD=0.0576p
+ PS=1.34u PD=0.74u
M$46 \$18 \$17 \$35 \$48 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.0576p
+ PS=0.74u PD=0.74u
M$47 \$35 \$17 \$18 \$48 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.0576p
+ PS=0.74u PD=0.74u
M$48 \$18 \$17 \$35 \$48 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.1026p
+ PS=0.74u PD=1.34u
M$49 \$36 \$18 \$19 \$49 sg13_lv_pmos L=0.13u W=0.18u AS=0.1026p AD=0.0576p
+ PS=1.34u PD=0.74u
M$50 \$19 \$18 \$36 \$49 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.0576p
+ PS=0.74u PD=0.74u
M$51 \$36 \$18 \$19 \$49 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.0576p
+ PS=0.74u PD=0.74u
M$52 \$19 \$18 \$36 \$49 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.1026p
+ PS=0.74u PD=1.34u
M$53 \$37 \$19 \$20 \$46 sg13_lv_pmos L=0.13u W=0.18u AS=0.1026p AD=0.0576p
+ PS=1.34u PD=0.74u
M$54 \$20 \$19 \$37 \$46 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.0576p
+ PS=0.74u PD=0.74u
M$55 \$37 \$19 \$20 \$46 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.0576p
+ PS=0.74u PD=0.74u
M$56 \$20 \$19 \$37 \$46 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.1026p
+ PS=0.74u PD=1.34u
M$57 \$66 \$4 \$65 \$68 sg13_lv_pmos L=0.13u W=0.155u AS=0.10085p AD=0.05585p
+ PS=1.34u PD=0.74u
M$58 \$65 \$4 \$64 \$68 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.05585p
+ PS=0.74u PD=0.74u
M$59 \$64 \$4 \$63 \$68 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.05585p
+ PS=0.74u PD=0.74u
M$60 \$63 \$4 \$67 \$68 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.10085p
+ PS=0.74u PD=1.34u
M$61 \$69 \$4 \$73 \$74 sg13_lv_pmos L=0.13u W=0.155u AS=0.10085p AD=0.05585p
+ PS=1.34u PD=0.74u
M$62 \$73 \$4 \$72 \$74 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.05585p
+ PS=0.74u PD=0.74u
M$63 \$72 \$4 \$71 \$74 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.05585p
+ PS=0.74u PD=0.74u
M$64 \$71 \$4 \$70 \$74 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.10085p
+ PS=0.74u PD=1.34u
M$65 \$78 \$4 \$77 \$79 sg13_lv_pmos L=0.13u W=0.155u AS=0.10085p AD=0.05585p
+ PS=1.34u PD=0.74u
M$66 \$77 \$4 \$76 \$79 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.05585p
+ PS=0.74u PD=0.74u
M$67 \$76 \$4 \$75 \$79 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.05585p
+ PS=0.74u PD=0.74u
M$68 \$75 \$4 \$80 \$79 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.10085p
+ PS=0.74u PD=1.34u
M$69 \$82 \$4 \$81 \$86 sg13_lv_pmos L=0.13u W=0.155u AS=0.10085p AD=0.05585p
+ PS=1.34u PD=0.74u
M$70 \$81 \$4 \$85 \$86 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.05585p
+ PS=0.74u PD=0.74u
M$71 \$85 \$4 \$84 \$86 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.05585p
+ PS=0.74u PD=0.74u
M$72 \$84 \$4 \$83 \$86 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.10085p
+ PS=0.74u PD=1.34u
M$73 \$87 \$4 \$90 \$92 sg13_lv_pmos L=0.13u W=0.155u AS=0.10085p AD=0.05585p
+ PS=1.34u PD=0.74u
M$74 \$90 \$4 \$91 \$92 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.05585p
+ PS=0.74u PD=0.74u
M$75 \$91 \$4 \$89 \$92 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.05585p
+ PS=0.74u PD=0.74u
M$76 \$89 \$4 \$88 \$92 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.10085p
+ PS=0.74u PD=1.34u
M$77 \$50 \$20 \$2 \$44 sg13_lv_pmos L=0.13u W=0.18u AS=0.1026p AD=0.0576p
+ PS=1.34u PD=0.74u
M$78 \$2 \$20 \$50 \$44 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.0576p
+ PS=0.74u PD=0.74u
M$79 \$50 \$20 \$2 \$44 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.0576p
+ PS=0.74u PD=0.74u
M$80 \$2 \$20 \$50 \$44 sg13_lv_pmos L=0.13u W=0.18u AS=0.0576p AD=0.1026p
+ PS=0.74u PD=1.34u
M$81 \$59 \$4 \$57 \$62 sg13_lv_pmos L=0.13u W=0.155u AS=0.10085p AD=0.05585p
+ PS=1.34u PD=0.74u
M$82 \$57 \$4 \$56 \$62 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.05585p
+ PS=0.74u PD=0.74u
M$83 \$56 \$4 \$60 \$62 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.05585p
+ PS=0.74u PD=0.74u
M$84 \$60 \$4 \$61 \$62 sg13_lv_pmos L=0.13u W=0.155u AS=0.05585p AD=0.10085p
+ PS=0.74u PD=1.34u
.ENDS VCO
