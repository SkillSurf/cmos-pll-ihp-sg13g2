* Extracted by KLayout with SG13G2 LVS runset on : 11/06/2025 07:50

.SUBCKT t2_freq_divider
X$1 \$4 \$1 \$28 t2_tie
X$2 \$1 \$4 \$6 \$14 \$5 \$16 \$19 t2_or4
X$3 \$4 \$1 \$26 t2_tie
X$8 \$1 \$4 \$26 \$30 \$30 \$5 \$32 t2_dff
X$9 \$4 \$20 \$11 \$1 \$7 t2_nand2
X$10 \$1 \$4 \$5 \$I40 \$I41 \$7 \$I39 t2_dff
X$11 \$1 \$9 \$4 \$3 \$I40 \$I39 t2_ha
X$12 \$1 \$4 \$12 \$I39 \$14 t2_xor2
X$13 \$1 \$4 \$5 \$I43 \$I44 \$7 \$I42 t2_dff
X$14 \$1 \$15 \$4 \$9 \$I43 \$I42 t2_ha
X$15 \$1 \$4 \$24 \$I42 \$16 t2_xor2
X$16 \$1 \$4 \$5 \$I46 \$I47 \$7 \$I45 t2_dff
X$17 \$1 \$28 \$4 \$15 \$I46 \$I45 t2_ha
X$18 \$1 \$4 \$33 \$I45 \$19 t2_xor2
X$19 \$1 \$4 \$5 \$I49 \$I50 \$7 \$I48 t2_dff
X$20 \$1 \$3 \$4 \$I20 \$I49 \$I48 t2_ha
X$21 \$1 \$4 \$8 \$I48 \$6 t2_xor2
.ENDS t2_freq_divider

.SUBCKT t2_or4 \$1 \$2 \$5 \$6 \$9 \$10 \$11
X$1 \$1 \$2 \$10 \$11 \$13 t2_or2
X$2 \$1 \$2 \$5 \$6 \$7 t2_or2
X$3 \$1 \$2 \$7 \$13 \$9 t2_or2
.ENDS t2_or4

.SUBCKT t2_tie \$1 \$4 \$5
M$1 \$6 \$3 \$4 \$4 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
M$2 \$4 \$2 \$2 \$4 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
M$3 \$1 \$3 \$3 \$1 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
M$4 \$5 \$2 \$1 \$1 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
.ENDS t2_tie

.SUBCKT t2_ha \$1 \$3 \$4 \$6 \$8 \$13
X$1 \$1 \$4 \$3 \$13 \$6 t2_and2
X$2 \$1 \$4 \$3 \$13 \$8 t2_xor2
.ENDS t2_ha

.SUBCKT t2_dff \$1 \$2 \$4 \$6 \$9 \$10 \$12
X$1 \$1 \$11 \$7 \$8 \$5 \$2 t2_nand3
X$2 \$2 \$1 \$10 \$8 t2_inverter
X$3 \$1 \$13 \$11 \$8 \$4 \$2 t2_nand3
X$4 \$1 \$12 \$9 \$7 \$4 \$2 t2_nand3
X$5 \$1 \$7 \$5 \$6 \$4 \$2 t2_nand3
X$6 \$2 \$11 \$9 \$1 \$12 t2_nand2
X$7 \$2 \$5 \$11 \$1 \$13 t2_nand2
.ENDS t2_dff

.SUBCKT t2_or2 \$1 \$2 \$4 \$5 \$9
X$1 \$2 \$5 \$5 \$1 \$8 t2_nand2
X$2 \$2 \$4 \$4 \$1 \$7 t2_nand2
X$3 \$2 \$8 \$7 \$1 \$9 t2_nand2
.ENDS t2_or2

.SUBCKT t2_and2 \$1 \$2 \$4 \$5 \$8
X$1 \$2 \$5 \$4 \$1 \$7 t2_nand2
X$2 \$2 \$7 \$7 \$1 \$8 t2_nand2
.ENDS t2_and2

.SUBCKT t2_inverter \$1 \$2 \$3 \$4
M$1 \$2 \$3 \$4 \$2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
M$2 \$1 \$3 \$4 \$1 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
.ENDS t2_inverter

.SUBCKT t2_nand3 \$1 \$2 \$3 \$4 \$5 \$12
M$1 \$3 \$2 \$6 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$2 \$6 \$4 \$10 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p
+ PS=0.74u PD=0.74u
M$3 \$10 \$5 \$1 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p
+ PS=0.74u PD=1.34u
M$4 \$12 \$2 \$3 \$12 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u
+ PD=0.68u
M$5 \$3 \$4 \$12 \$12 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.057p PS=0.68u
+ PD=0.68u
M$6 \$12 \$5 \$3 \$12 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u
+ PD=1.28u
.ENDS t2_nand3

.SUBCKT t2_xor2 \$1 \$2 \$4 \$5 \$11
X$1 \$2 \$5 \$4 \$1 \$6 t2_nand2
X$2 \$2 \$9 \$10 \$1 \$11 t2_nand2
X$3 \$2 \$5 \$6 \$1 \$9 t2_nand2
X$4 \$2 \$6 \$4 \$1 \$10 t2_nand2
.ENDS t2_xor2

.SUBCKT t2_nand2 \$1 \$2 \$3 \$4 \$5
M$1 \$4 \$2 \$6 \$4 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$2 \$6 \$3 \$5 \$4 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$3 \$1 \$2 \$5 \$1 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u
+ PD=0.68u
M$4 \$5 \$3 \$1 \$1 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u
+ PD=1.28u
.ENDS t2_nand2
