** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_ha_tb.sch
**.subckt t2_ha_tb
x1 VDD GND A B S C t2_ha
VinA A GND dc 0 ac 0 pulse(0, 1.2, 0, 50p, 50p, 1.25n, 2.5n)
VinB B GND dc 0 ac 0 pulse(0, 1.2, 0, 50p, 50p, 2.5n, 5n)
Vs VDD GND 1.2
* noconn S
* noconn C
**** begin user architecture code


.param temp=27
.control
save all
tran 10p 10n
write tran_t2_ha.raw
.endc



.lib cornerMOSlv.lib mos_ff

**** end user architecture code
**.ends

* expanding   symbol:  t2_ha.sym # of pins=6
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_ha.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_ha.sch
.subckt t2_ha VDD VSS inA inB sum cout
*.iopin VSS
*.ipin inA
*.ipin inB
*.opin sum
*.iopin VDD
*.opin cout
x1 VDD VSS inA inB sum t2_xor2
x2 VDD VSS inA cout inB t2_and2
.ends


* expanding   symbol:  t2_xor2.sym # of pins=5
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_xor2.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_xor2.sch
.subckt t2_xor2 VDD VSS inA inB out
*.iopin VSS
*.ipin inA
*.ipin inB
*.opin out
*.iopin VDD
x1 VDD inA inB net1 VSS t2_nand2
x2 VDD inA net1 net3 VSS t2_nand2
x3 VDD net1 inB net2 VSS t2_nand2
x4 VDD net3 net2 out VSS t2_nand2
.ends


* expanding   symbol:  t2_and2.sym # of pins=5
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_and2.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_and2.sch
.subckt t2_and2 VDD VSS inA out inB
*.iopin VSS
*.ipin inA
*.ipin inB
*.opin out
*.iopin VDD
x1 VDD inA inB net1 VSS t2_nand2
x2 VDD net1 net1 out VSS t2_nand2
.ends


* expanding   symbol:  t2_nand2.sym # of pins=5
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand2.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_nand2.sch
.subckt t2_nand2 VDD inA inB out VSS
*.iopin VSS
*.ipin inA
*.ipin inB
*.opin out
*.iopin VDD
XM1 out inA VDD VDD sg13_lv_pmos w=0.3u l=0.15u ng=1 m=1
XM2 out inB VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
XM3 out inB net1 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM4 net1 inA VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
