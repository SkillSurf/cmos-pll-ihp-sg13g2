** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/11Stage_vco_new.sch
.subckt 11Stage_vco_new VPWR VGND vctl Vout
*.PININFO VPWR:B VGND:B vctl:I Vout:O
M21 mirror_pg mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
M22 net1 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
M23 net2 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
M24 net3 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
M25 mirror_pg vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
M26 net9 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
M28 net7 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
M29 net13 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
M30 net12 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
M31 net10 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
M32 net11 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
M33 net15 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
M34 net16 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
M35 net20 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
M36 net19 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
M37 net24 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
M38 net23 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
M39 net21 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
M40 net22 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
M41 net31 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
M42 net30 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
M43 net28 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
M44 net29 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
M1 net8 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
C12 VGND net4 cap_cmim w=6.99e-6 l=6.99e-6 m=1
C1 VGND net5 cap_cmim w=6.99e-6 l=6.99e-6 m=1
C2 VGND net6 cap_cmim w=6.99e-6 l=6.99e-6 m=1
C3 VGND net14 cap_cmim w=6.99e-6 l=6.99e-6 m=1
C4 VGND net26 cap_cmim w=6.99e-6 l=6.99e-6 m=1
C5 VGND net17 cap_cmim w=6.99e-6 l=6.99e-6 m=1
C6 VGND net18 cap_cmim w=6.99e-6 l=6.99e-6 m=1
C7 VGND net25 cap_cmim w=6.99e-6 l=6.99e-6 m=1
C8 VGND net27 cap_cmim w=6.99e-6 l=6.99e-6 m=1
C9 VGND net32 cap_cmim w=6.99e-6 l=6.99e-6 m=1
C10 VGND feedback cap_cmim w=6.99e-6 l=6.99e-6 m=1
C11 VGND Vout cap_cmim w=6.99e-6 l=6.99e-6 m=2
x13 net1 VPWR feedback net4 VGND net9 vco_inverter
x1 net2 VPWR net4 net5 VGND net8 vco_inverter
x2 net3 VPWR net5 net6 VGND net7 vco_inverter
x3 net13 VPWR net6 net14 VGND net10 vco_inverter
x4 net12 VPWR net14 net26 VGND net11 vco_inverter
x5 net15 VPWR net26 net17 VGND net20 vco_inverter
x6 net16 VPWR net17 net18 VGND net19 vco_inverter
x7 net24 VPWR net18 net25 VGND net21 vco_inverter
x8 net23 VPWR net25 net27 VGND net22 vco_inverter
x9 net31 VPWR net27 net32 VGND net28 vco_inverter
x10 net30 VPWR net32 feedback VGND net29 vco_inverter
x11 VPWR VPWR feedback Vout VGND VGND vco_inverter
.ends

* expanding   symbol:  vco_inverter.sym # of pins=6
** sym_path: /foss/designs/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/vco_inverter.sym
** sch_path: /foss/designs/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/vco_inverter.sch
.subckt vco_inverter VPWR VPB A Y VNB VGND
*.PININFO VPWR:B VGND:B A:I Y:O VPB:B VNB:B
M2 Y A VPWR VPB sg13_lv_pmos w=2u l=0.13u ng=1 m=1
M1 Y A VGND VNB sg13_lv_nmos w=1u l=0.13u ng=1 m=1
.ends

