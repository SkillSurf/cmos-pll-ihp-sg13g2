** sch_path: /foss/designs/Team1/PLL_Completed/PLL_Completed_tb.sch
**.subckt PLL_Completed_tb
x1 Fref UP net1 DN net2 Ffeed PFD
x2 Vdd ICP GND net1 UP VCON net2 DN CP_LF
x3 Vdd VCO_OUT VCON GND VCO_3Stages
x4 Vdd Ffeed VCO_OUT GND Div8F
V1 Vdd GND 1.2
I0 Vdd ICP 80u
Vin1 Fref GND dc 0 ac 0 pulse(0, 1.2, 0, 10p, 10p, 2.5n, 5n)
**** begin user architecture code


.param temp=27
.control
save all
.options maxstep=10n reltol=1e-3 abstol=1e-6
tran 50p 600n
plot v(Fref)+10 v(Ffeed)+8 v(UP)+6 v(DN)+4 v(VCO_OUT)+2 v(VCON) xlimit 400n 600n
fft v(VCO_OUT)
plot db(mag(v(VCO_OUT))) xlabel 'Frequency ' xlimit 0 2Gig
.endc


 .lib cornerMOSlv.lib mos_tt

**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/Team1/PFD/PFD.sym # of pins=6
** sym_path: /foss/designs/Team1/PFD/PFD.sym
** sch_path: /foss/designs/Team1/PFD/PFD.sch
.subckt PFD Fref UP UPB DN DNB Ffeed
*.ipin Fref
*.ipin Ffeed
*.opin UP
*.opin UPB
*.opin DN
*.opin DNB
x1 Fref net1 Fref 2NAND
x2 UPB net3 net1 2NAND
x3 net3 net5 net4 2NAND
x4 net5 net4 net6 2NAND
x5 net6 net7 net8 2NAND
x6 Ffeed net2 Ffeed 2NAND
x7 net2 net9 DNB 2NAND
x8 net7 net8 net9 2NAND
x9 net8 net11 net9 2NAND
x10 net3 net10 net5 2NAND
x11 net10 net12 net10 2NAND
x12 net11 net13 net11 2NAND
x13 net12 net6 net13 2NAND
x14 UPB UP UPB 2NAND
x15 DNB DN DNB 2NAND
x16 UPB net3 net5 net6 3NAND
x17 DNB net6 net8 net9 3NAND
.ends


* expanding   symbol:  /foss/designs/Team1/CP_LF/CP_LF.sym # of pins=8
** sym_path: /foss/designs/Team1/CP_LF/CP_LF.sym
** sch_path: /foss/designs/Team1/CP_LF/CP_LF.sch
.subckt CP_LF VDD ICP VSS UPB UP VCON DNB DN
*.iopin VDD
*.iopin ICP
*.iopin VSS
*.ipin UPB
*.ipin UP
*.ipin DNB
*.ipin DN
*.opin VCON
XM1 net1 net1 VDD VDD sg13_lv_pmos w=0.5u l=0.2u ng=1 m=1
XM2 net4 net1 VDD VDD sg13_lv_pmos w=0.5u l=0.2u ng=1 m=1
XM3 net3 net4 VDD VDD sg13_lv_pmos w=1.1u l=0.2u ng=1 m=10
XM4 net4 ICP net3 VDD sg13_lv_pmos w=1.1u l=0.2u ng=1 m=10
XM5 ICP ICP VDD VDD sg13_lv_pmos w=4u l=0.5u ng=1 m=1
XM6 net5 net4 VDD VDD sg13_lv_pmos w=1.1u l=0.2u ng=1 m=10
XM7 VCON ICP net5 VDD sg13_lv_pmos w=1.1u l=0.2u ng=1 m=10
XM8 net6 net6 VDD VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=10
XM9 net8 net6 VDD VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=10
XM10 ICP ICP VSS VSS sg13_lv_nmos w=2u l=0.2u ng=1 m=1
XM11 net4 UP net2 VSS sg13_lv_nmos w=2u l=0.13u ng=1 m=1
XM12 net1 UPB net2 VSS sg13_lv_nmos w=2u l=0.13u ng=1 m=1
XM13 net2 ICP VSS VSS sg13_lv_nmos w=2u l=0.2u ng=1 m=1
XM14 net8 DNB net7 VSS sg13_lv_nmos w=2u l=0.13u ng=1 m=1
XM15 net6 DN net7 VSS sg13_lv_nmos w=2u l=0.13u ng=1 m=1
XM16 net7 ICP VSS VSS sg13_lv_nmos w=2u l=0.2u ng=1 m=1
XM19 VCON ICP net10 VSS sg13_lv_nmos w=10u l=0.2u ng=1 m=1
XM20 net10 net8 VSS VSS sg13_lv_nmos w=10u l=0.2u ng=1 m=1
XM21 net8 ICP net9 VSS sg13_lv_nmos w=10u l=0.2u ng=1 m=1
XM22 net9 net8 VSS VSS sg13_lv_nmos w=10u l=0.2u ng=1 m=1
R1 VCON net11 1k m=1
C1 net11 VSS 50f m=1
C2 VCON VSS 10f m=1
XM23 ICP ICP VSS VSS sg13_lv_nmos w=2u l=0.2u ng=1 m=1
.ends


* expanding   symbol:  /foss/designs/Team1/VCO/VCO_3Stages.sym # of pins=4
** sym_path: /foss/designs/Team1/VCO/VCO_3Stages.sym
** sch_path: /foss/designs/Team1/VCO/VCO_3Stages.sch
.subckt VCO_3Stages VDD VOUT VCON VSS
*.iopin VDD
*.iopin VSS
*.ipin VCON
*.opin VOUT
XM1 net1 net1 VDD VDD sg13_lv_pmos w=3u l=0.13u ng=1 m=1
XM2 net9 net1 VDD VDD sg13_lv_pmos w=3u l=0.13u ng=1 m=1
XM3 net8 net1 VDD VDD sg13_lv_pmos w=3u l=0.13u ng=1 m=1
XM4 net6 net1 VDD VDD sg13_lv_pmos w=3u l=0.13u ng=1 m=1
XM5 net1 VCON VSS VSS sg13_lv_nmos w=2u l=0.13u ng=1 m=1
XM6 net10 VCON VSS VSS sg13_lv_nmos w=2u l=0.13u ng=1 m=1
XM7 net7 VCON VSS VSS sg13_lv_nmos w=2u l=0.13u ng=1 m=1
XM8 net5 VCON VSS VSS sg13_lv_nmos w=2u l=0.13u ng=1 m=1
C2 VOUT VSS 10f m=1
x1 net9 net10 net2 net4 net2 New_2NAND
x2 net8 net7 net4 net3 net4 New_2NAND
x3 net6 net5 net3 net2 net3 New_2NAND
x4 VDD VSS net2 VOUT net2 New_2NAND
.ends


* expanding   symbol:  /foss/designs/Team1/FD/Div8F/Div8F.sym # of pins=4
** sym_path: /foss/designs/Team1/FD/Div8F/Div8F.sym
** sch_path: /foss/designs/Team1/FD/Div8F/Div8F.sch
.subckt Div8F VDD FOUT FIN VSS
*.opin FOUT
*.ipin FIN
*.iopin VDD
*.iopin VSS
x1 VDD net2 net1 FIN net2 VSS DFlop
x2 VDD net4 net3 net1 net4 VSS DFlop
x3 VDD net5 FOUT net3 net5 VSS DFlop
.ends


* expanding   symbol:  /foss/designs/Team1/2NAND/2NAND.sym # of pins=3
** sym_path: /foss/designs/Team1/2NAND/2NAND.sym
** sch_path: /foss/designs/Team1/2NAND/2NAND.sch
.subckt 2NAND A Y B
*.ipin B
*.opin Y
*.ipin A
XM1 Y A net1 net1 sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM2 Y B net1 net1 sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM3 Y B net2 GND sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM4 net2 A GND GND sg13_lv_nmos w=1u l=0.13u ng=1 m=1
V1 net1 GND 1.2
.ends


* expanding   symbol:  /foss/designs/Team1/3NAND/3NAND.sym # of pins=4
** sym_path: /foss/designs/Team1/3NAND/3NAND.sym
** sch_path: /foss/designs/Team1/3NAND/3NAND.sch
.subckt 3NAND Y A B C
*.ipin A
*.ipin B
*.ipin C
*.opin Y
XM1 Y A Vdd Vdd sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM2 Y B Vdd Vdd sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM3 Y C Vdd Vdd sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM4 Y A net1 GND sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM5 net1 B net2 GND sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM6 net2 C GND GND sg13_lv_nmos w=1u l=0.13u ng=1 m=1
V1 Vdd GND 1.2
.ends


* expanding   symbol:  /foss/designs/Team1/New_2NAND/New_2NAND.sym # of pins=5
** sym_path: /foss/designs/Team1/New_2NAND/New_2NAND.sym
** sch_path: /foss/designs/Team1/New_2NAND/New_2NAND.sch
.subckt New_2NAND VDD VSS A Y B
*.ipin B
*.opin Y
*.ipin A
*.iopin VDD
*.iopin VSS
XM1 Y A VDD VDD sg13_lv_pmos w=3u l=0.13u ng=1 m=1
XM2 Y B VDD VDD sg13_lv_pmos w=3u l=0.13u ng=1 m=1
XM3 Y B net1 VSS sg13_lv_nmos w=2u l=0.13u ng=1 m=1
XM4 net1 A VSS VSS sg13_lv_nmos w=2u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  /foss/designs/Team1/DFlop/DFlop.sym # of pins=6
** sym_path: /foss/designs/Team1/DFlop/DFlop.sym
** sch_path: /foss/designs/Team1/DFlop/DFlop.sch
.subckt DFlop VDD D Q CLK QBAR VSS
*.iopin VDD
*.iopin VSS
*.ipin D
*.ipin CLK
*.opin Q
*.opin QBAR
XM1 net1 D VDD VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM2 net4 CLK VDD VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM3 QBAR net4 VDD VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM4 Q QBAR VDD VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM5 net2 CLK net1 VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM6 QBAR CLK net5 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM7 net4 net2 net3 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM8 net2 D VSS VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM9 net3 CLK VSS VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM10 net5 net4 VSS VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM11 Q QBAR VSS VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
C1 QBAR VSS 10f m=1
C2 Q VSS 10f m=1
.ends

.GLOBAL GND
.end
