** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/dff_nclk_tb.sch

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.include /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice

**.subckt dff_nclk_tb
Vdin D GND dc 0 ac 0 pulse(0, 1.2, 0, 100p, 100p, 12.5n, 25n)
Vclk nCLK GND dc 0 ac 0 pulse(0, 1.2, 0, 100p, 100p, 6.25n, 12.5n)
Vrst nRST GND dc 0 ac 0 pulse(0, 1.2, 0, 100p, 100p, 40n, 75n)
* noconn nQ
* noconn Q
x1 nCLK Q D nQ nRST net1 GND dff_nclk
Vs net1 GND 1.2
**** begin user architecture code


.param temp=27
vvdd vdd 0 dc 1.2
vvss vss 0 0
.control
pre_osdi ./psp103_nqs.osdi
save all
tran 50p 75n

write tran_dff_nclk.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  dff_nclk.sym # of pins=7
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/dff_nclk.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/dff_nclk.sch
.subckt dff_nclk nCLK Q D nQ nRST VDD VSS
*.ipin nCLK
*.ipin D
*.ipin nRST
*.opin Q
*.opin nQ
*.iopin VSS
*.iopin VDD
x1 net1 D Q nQ nRST VDD VSS sg13g2_dfrbp_1
x2 nCLK VDD VSS net1 sg13g2_inv_1
.ends

.GLOBAL GND
.end
