** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Team 2 Design/design_data/xschem/t2_inverter.sch
.subckt t2_inverter VP A Y VN
*.PININFO VP:B VN:B A:I Y:O
M2 Y A VP VP sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M1 Y A VN VN sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends
