** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/dff_tb.sch

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.include /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice

**.subckt dff_tb
x1 clk d q qn net1 VDD VSS sg13g2_dfrbp_1
Vclk clk GND dc 0 ac 0 pulse(0, 1.2, 6.25n, 100p, 100p, 6.25n, 12.5n)
Vdin d GND dc 0 ac 0 pulse(0, 1.2, 0, 100p, 100p, 12.5n, 25n)
* noconn q
* noconn qn
Vrst net1 GND dc 0 ac 0 pulse(0, 1.2, 0, 100p, 100p, 40n, 75n)
**** begin user architecture code


.param temp=27
vvdd vdd 0 dc 1.2
vvss vss 0 0
.control
pre_osdi ./psp103_nqs.osdi
save all
tran 50p 75n

write tran_dff.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
