** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/2-bit_freq_divider_tb.sch

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.include /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice

**.subckt 2-bit_freq_divider_tb
Vs VDD GND 1.2
Vclk CLK_IN GND dc 0 ac 0 pulse(0, 1.2, 0, 100p, 100p, 6.25n, 12.5n)
* noconn CLK_OUT
Ven EN GND dc {EN}
Va0 A0 GND dc {A0}
Va1 A1 GND dc {A1}
x1 VDD GND A0 CLK_OUT CLK_IN EN A1 2-bit_freq_divider
**** begin user architecture code


.meas tran tperiod_in TRIG v(clk_in) VAL=0.5 FALL=1 TARG v(clk_in) VAL=0.5 FALL=2
.meas tran freq_in PARAM = '1e-6/tperiod_in'

.meas tran tperiod_out TRIG v(clk_out) VAL=0.5 FALL=1 TARG v(clk_out) VAL=0.5 FALL=2
.meas tran freq_out PARAM = '1e-6/tperiod_out'

.meas tran tdelay TRIG v(clk_in) VAL=0.5 RISE=1 TARG v(clk_out) VAL=0.5 RISE=1




.param EN = 1.2

.param A0 = 1.2
.param A1 = 1.2




.param temp=27

.control
pre_osdi ./psp103_nqs.osdi
save all
tran 50p 150n

write tran_2-bit_freq_divider.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  2-bit_freq_divider.sym # of pins=7
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/2-bit_freq_divider.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/2-bit_freq_divider.sch
.subckt 2-bit_freq_divider VDD VSS A0 CLK_OUT CLK_IN EN A1
*.ipin CLK_IN
*.ipin EN
*.ipin A0
*.ipin A1
*.opin CLK_OUT
*.iopin VSS
*.iopin VDD
x1 VDD GND nEQ0 net1 CLK net2 DIV_RST A0 freq_div_cell
x2 VDD GND nEQ1 net2 CLK Cout DIV_RST A1 freq_div_cell
x3 net1 VDD VSS sg13g2_tiehi
* noconn Cout
x4 nEQ0 nEQ1 VDD VSS DIV_RST sg13g2_or2_1
x5 DIV_RST CLK_OUT net3 net3 net4 VDD GND dff_nclk
x6 net4 VDD VSS sg13g2_tiehi
* noconn CLK_OUT
x7 CLK_IN EN VDD VSS CLK sg13g2_nand2_1
.ends


* expanding   symbol:  freq_div_cell.sym # of pins=8
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/freq_div_cell.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/freq_div_cell.sch
.subckt freq_div_cell VDD VSS DIV Cin CLK Cout nRST BIT
*.ipin Cin
*.ipin CLK
*.ipin nRST
*.ipin BIT
*.opin DIV
*.opin Cout
*.iopin VSS
*.iopin VDD
x1 net2 net1 Cin VDD VSS Cout half_add
x2 CLK net2 net1 net3 nRST VDD VSS dff_nclk
x3 net2 BIT VDD VSS DIV sg13g2_xor2_1
* noconn #net3
.ends


* expanding   symbol:  dff_nclk.sym # of pins=7
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/dff_nclk.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/dff_nclk.sch
.subckt dff_nclk nCLK Q D nQ nRST VDD VSS
*.ipin nCLK
*.ipin D
*.ipin nRST
*.opin Q
*.opin nQ
*.iopin VSS
*.iopin VDD
x1 net1 D Q nQ nRST VDD VSS sg13g2_dfrbp_1
x2 nCLK VDD VSS net1 sg13g2_inv_1
.ends


* expanding   symbol:  half_add.sym # of pins=6
** sym_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/half_add.sym
** sch_path: /foss/designs/PROJECTS/cmos-pll-ihp-sg13g2/Combined Design/design_data/xschem/half_add.sch
.subckt half_add inA sum inB VDD VSS cout
*.ipin inA
*.ipin inB
*.opin sum
*.opin cout
*.iopin VSS
*.iopin VDD
x1 inA inB VDD VSS sum sg13g2_xor2_1
x2 inA inB VDD VSS cout sg13g2_and2_1
.ends

.GLOBAL GND
.end
