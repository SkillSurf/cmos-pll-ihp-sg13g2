** sch_path: /foss/designs/Team1/New_2NAND/New_2NAND_tb.sch
**.subckt New_2NAND_tb Vout
*.opin Vout
Vin VB GND dc 0 ac 0 pulse(0, 1.2, 0, 10p, 10p, 2n, 4n)
Vin1 VA GND dc 0 ac 0 pulse(0, 1.2, 5n, 10p, 10p, 3n, 6n)
C1 Vout GND 100f m=1
V1 net1 GND 1.8
x1 net1 GND VA Vout VB New_2NAND
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt



.param temp=27
.control
save all
tran 1n 20n
plot v(VA)+4 v(VB)+2 v(Vout)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/Team1/New_2NAND/New_2NAND.sym # of pins=5
** sym_path: /foss/designs/Team1/New_2NAND/New_2NAND.sym
** sch_path: /foss/designs/Team1/New_2NAND/New_2NAND.sch
.subckt New_2NAND VDD VSS A Y B
*.ipin B
*.opin Y
*.ipin A
*.iopin VDD
*.iopin VSS
XM1 Y A VDD VDD sg13_lv_pmos w=3u l=0.13u ng=1 m=1
XM2 Y B VDD VDD sg13_lv_pmos w=3u l=0.13u ng=1 m=1
XM3 Y B net1 VSS sg13_lv_nmos w=2u l=0.13u ng=1 m=1
XM4 net1 A VSS VSS sg13_lv_nmos w=2u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
